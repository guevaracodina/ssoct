��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ��p"���C��T�fX��k�+��)��6�'�3��$���)��2�+�
�#�7��Ib����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�o ���`=<��3+�)L�Q*$�:-m��]x[;_ߐ��c�L2��0��z�����9� �?Q����ھO��� �ߣNA�B�1"���;3}��=�g��N��D.݁z�.<�f�ӁD�x}��u=k+��	���F�k_	����~T���nۘ_���Ѩ���^S�z��ۅ��Ѩ{Jf�D9:k(��ѻ](� |A�B�F��:��$/�}֏��!�i��q��&)��;��>\���O��r���Y��N�j�㐫WW��C��/C2�>��;�;�?�H�QI��CR�1l�զ�N����NLE�J'�m��W1�l|�9H]B���#ű��l�j��Z[e��=@굁�,���D�=�'��>���|�VUg!�A�6�m�x�F*>�i�#�~���0�=�M��]s�������bI�� �.�fdB09$H� \u�-�8�z�Ğa�Lr�-P�MH�,e��0��p�����A��$6��$��Z6����,33��'��h����kY��X��/�p� 
?���懣X�G���Z��X��{����� j�`-�Ti4�'JH�(���V��/B�8���ZـS��P�r��a>q8V����Q���-�/G��^�`:V��Q��1*��!���CL��	X�F3�OYۓ�EB&y�A�	��Ӡ�mA|B�Cu�ٵ����7���C��Y�o�:���)�n��D�2�TJW`���/k�b�k[B>Ǖ��r�N\���94Q}F6��#�Ԉ��81.ƕ�������!�:)șIS�#"_�#L�`ƍnA�^�<�>C�
��\b�� �T��	-�Kqt�ey3�x�b�0#�gR�&�@��(��|��J����fr�o�#�D�#uD(x�?�9E��]��Z��`����(f�ܲ�*�-��H��!X��D:t��3 䇏2pVw�r]��"{YJf���x�� �{*��Ɏ�񮤀Q��%u�ݶ
�3|LOe�Z)ZS%�"�lhc_ID��)[#�sL>�B>K�iH	�y3��	�yňr�+1B��z��[�Bf)�er9����H�Z��\�:�Y��G�ʈ�?AȤ8�:�M^5�CU�zn&��J��䎕L~�W<K��[z��x��7�g����6�"���c�n7�z���C��^e��e�l�&Q�9nkI��4�S��ϵT#�[PzD���J�󒙐�2���F��Y�QX0TL^�Lvgx<�u}5oh�aʜ����������XZ��
)1��(3�($	����ĂA����K:T�8�syeTs���$���uQ��ӈ�*�n)xkЦ��?}q߹Q�G.Jl�~�=E��X��^"�����ym9I��fZ��	50���y=6���^���vD��z�`�j/��q�.��Ǳ1Z��|����Q'W6�Gu��U��ί�%0��ՙ��S�8�O��o��r"^	�#��oi�w�J��h����k�;?9���]��(��6���%�&��+L��R�>K[N<a0�8U���rۯ��%F�*�]"K
�q�"J@!a�d��͙�fJ��L��f���;�ΗK�JU�x>��6��u��sh7-��5k�IU�_g��_�;�~�mO��W~��i��L��u�"	
�./�Qڗ��ת`�q��蛡S�����ƹH��|X�0�/���9�x�r��
�>Șh����s�]���M;�	��/�C�Su�	�.����� Y��S�.��=��	��c�Iת�t�����6��?��d��:-ph+DZ/������IpO�Ƹ�F*�^#X�44�D�U��hXE���V*��Uնg��� �����̃)�m���l������r�*u�^��T�/d�*RB�Q�/��h��B!9�W�qg�2�&E>՗����ak�L��lw�?�����H橘$zB�����7�H��I�
���؛J�V�&,�6z�'�� �����Q+b5l#&Zg�� c�,o=G�ޓ���K�2���*����&�J8)�HMG��OV���D�2�re͕L��N`Ǧ��A�^���g{(!Υ�غ~t��S�JHO@�<���zV���J��X��K^p�z钌���)����'��s2ǉ*�f�D�B.%%�b��Z(z�s$��S�֖�$�4O�i9I��(k�f���OB��a���55�Z��>�d�z#9�e�?�����Q37��[�?^D_�.��\�J��B_�~��u�O*���1L��A݌��m�s?�(̻T��|��`���v.� @%S���f��U��Qp�J+�תJ����`�=w����9}n�L������+1�qB�{��?���.�Px6'�j�jS(��C���/B��S'����Ȋ�!�X��\X428�8�e>J�VT{�m��|zX3�|����%��_O�YW�ѠT.Y9��uB7w�
�����ݷl�a��)]�� թ=pT��k��}�\O+�Hu�U,~��az������s���
�<��|�A6I��9B��6 o�(�\.U���P�!u[<RU��\wo��Ox��1<g�>���C��䠠 CA���V7��T0f�)��Ĝ�EKR�.����*��(���:�Z�ږ�zM#�:�[�������P9�qZ��p4o�͊6��IWb��*=8�O{����UN�.�����R�B8�^�dӕ^�3-%k{	� :��c3�co����s�U�G��yəm``�H԰)�$���d�e��X�L���7��H.��g��cf���IT�Qm=�o�e� ���O�T�������k�͙�	H ����=��	�h�v�"�c%/,s���Mvc*/�q�v}-�P���j2�1e͉�����/s�!�T���s �`z`|'���#�y�Ϯ���KMu�}����o��=�t��Z[8#�� �O�)9'����F;����YP-v���|���$}�q��2�QW�������ϯsgkY>w���s���Y!u$~������,9Bг@�JT���&"��32V�����xA�3k�$�z� *j����.E&VdF���F��Yr3/�`7��#��D�sI�|����tq�"�0by�c�{��W����p\Yx|_�7x'��{A��@�<b��6��k�O����4GK=�-M��;$2-pN�q��R==�=��