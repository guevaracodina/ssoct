��/  S����3�c�ub��_NЀP���t�,ï�!U;�P{�g��Oj*�x �*�'|�N�Q]/]X	�b4)�Ob��8�O��ȸ�O_�&��*��2����K�I:[�Q�Ar���C�T&���Ͽ.W�����C�e8�<K��L�J[�(M;���B;"|�!���6?����d�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P�!�t������CC����<{)]%e�Щ�K,��YV�ґ4s�^[	�8H1��â������M�4Z��5b��O��u5��g�Y?������uXe�A�'P$v�_ye?�܇�_�Y���YWv�x��kٻi.���}��Z0]"��63�.�dC�T���gb����:�]*�>��ޘ�xW�c�`d��/820�/J���ˏ�-X��!��	;�A��o�l�������(����(�(x'fef�+�W�cEKW@�n���XD�4������J�7
�}qV�Y��cc��g���C0S4��񭸖�?�&��j�~�7%��r#�~��B���a�]>��m�IOs�M�-�gm8����)�.R��eZ����8�>�J�?S�L�\ҔY�9ʷ��t���P<n˄�}�Y�Pw0��簘�5� ��I�KZ���bS��|mf�ޒ*C�{���wi��	O�!{9B�2}�'&ZC��nxw�J.4��f�������������D���G���Izф�mGq4ό��<���D�#�#lª��+ 
w�l�T�1�nJy�6h->�1����ʼA}98Ǣe�t;Zs���Z��A�(1-�IEW:���p�HP�}Q�%�Uk� Ut��+~�r%k�![q�+���JnU2o-2C�������y\��m��"������e���*зs.�~Iؖh��h$8(4�_���NN*.�BԀ�U'�������E����¦ʒ8�?D��\��6V��Qȟ����������u��[N�$s'\�Q��G",��O)�B�cؕSTd�@��[q��_�Ո�k��]�bO�Ct?_��^����W��x�?�8���e|����Z�c��Óv�����a�����I�V �,$�L�i��D�ԍ�v7�v�evUx������5��]Yd�'�~��t��t��I�n9��[q.��L�&�B�ZP�f�3�0Ԙ�%{i�	��F��s��j��]wI! �E���(h��J3�T���+*a�*�I�l��k򃐄������r0/��2����Ql��V��Lt�]�%��*Bʦ���vg4hB����*}Nki\ǴU���|��� H+5�KH�5d������\��7��95��]c~���8*M��h��NX/�ݺU��wǓ��;�a*��O�S��ǜ0�Jq���6㶖_��T���
��=x	&�epŪYa��x�|?aη�'m��#55�H�6�_�����V��eC��gE�\� /�Ԏ@�3�2�_����`\Z������̧��N�Le���G2}j���O/4,�=����~r2��E:v^�E���$S�n*a�����	�'�Y�V ��>��L"�u����wμ���U	Y� �M�(y��J�����d���;��ټ,�Gu'^�D`��� � ��ۈ�ݷD2�-��yN�d'K3Uc�ۨ:7k�č_�7��+�*����oS�N���������B�tk�ڪ)��ʂe����hS6���t%p����ֈ^�H�H�y?�R��k���2b^{*��AN@��68Ā��	�h0���u�T
������T�#���lt��_�z:���4I��O,�a���|pd��9�J�}���%�5�!,H�W�Zyr���T��F�g��z�h6��>C��Ge?�,��W��G8e�**���]n�C������N� 0Ά�����v֨BB�����:�5z��9��LsR�5`�� �T�`��ۧ��4��5~��e����G��ȣij;�?K�/�����~w)�&�u���hE��2��W� �{]���l�Ž;7Y�y4�xB�Z6bԻty�"�HJe8>���$�0}q�*�犇��,\��&/����C�uߖ��j��L䩊r�e ��k����x�E�iP�.��5F�JW;K-�T#� ��o{��\�IM���q�N}��������*�u�t�p��
��?�ւf�$��`�6ޮ���`�RY�5̽�`�պr"�L$�2 7e�Ah�зoT"~��[��C�K���a{�g�_>Ŋ N�R��`�.<]HC�4n7P<�$�B^�]����F:�J{�5eƓ%�q�K㝾U~d�Ԑ���o��v4��P�ZR�z����hl��7j�����
��Ԍ���1��������7��YG$�����Eᒻq�U4�8���7ZK>�<~���x���7dd}��]��FC��\edb|���b4��^�`�Z�s3=ix��=��g�	tS���0'�O�
����s�1����S<��
Hͻ���O�����Z\w%�>��7�ؤ�lu�>�ؕw 5���{DeLu'�r0�Ѝ��0�5��4bj�)��s�?r~�A���Yw� ]o�x�L�(�e=ƙFό�̳s=i-��m]]�.������պ�  xıCy3�Qi��]"Ϥ���g�Q��e�`���,B��\�����g�t�k���z�b�|��J��T�2׻�]����T�V�3��B 2�h����O �7���-ķ�Ю�F�F]Ӭ�u��΢[�^j��t��{�1�\�
�V���Z�"�NUO���\g2qh�pQ����|���Y�Ҭ�	��>9�I��V]y���Ņ��s�|VZˋd�����bBA���H0��@G��@��'��xZ��z3�B��,��e�c�ܱp��G$}��fyGtF��F>U��_���>�Kx$=4ꬸ��:14�KÒ�	����q���,�%��6�U� &�BH��!0�+�S��"B�(݃<��
�+ԝ۪�JS�HH�C�l�P����O,�.M	r�Պ�\bΑ<%��R�qv=�2�����E���_���]�uO ?���Ҷ��s�}���R�J�b����5#F� ���N6*݅>�+���uI¬�ȼ�����=Rڿ!��>03�G,�J$�#C��#�֔��R�Q��Q4]x%��9d�vŞ��څ�ߏ�?��7�N��..���Ů��;L�����='����1V|�TZh�i�ȟ��Kj�/E�\k�/ ����z�]_h��I���ʀN�j8��7�P=Y��c�0��������f�y� 	+��\U�RP"WgXcoG4���%13�0����K�`U-�m���Yշ�\$r3���p��n�)�j�T�n�5���[����94�����7��{�cd&�x��d\u�U@:�b��:��U4�Ú:
�"�c�U��M�ó�"���ͧ�D���E�W;h�	 �T���=�i},o�֜4���yW��W��A�BU���� NG� :<ݪ���64>�g**fg�ڍ�pn��T�؛ʣ-���w�ӡ��̂$`��&��T/�ϥ]�s�'Y1Z�U���m ����c<z��Ž-h7�x3	��_�7�A\p�Ć.Xrr�֮Q�Z��D9?�]zXԴk�Τ_�&�%�L ڦ�N`#��5�9d�����8Le�p#ڂfZ'5���w)_�Ґ@VkM�D�4ϫ%�BV*D���AAG��T�A�ͩ�#@Ewpxg
�	[�+�=�h?O��O��dV��S��@.�5��G��0�9)����B<;�f��+���I�X��p��@��&hUn�Y��y�h�lN7a4�b�g|��B���`5A�!
w�t���F�6F�Y	v᡺d���-@�gŷHt�)Q]2�PBMaj���	��ߓ����������9��1�@�D��d1�FsJH�Z��I1gЦ��ٳX< ��hd���@�����Q�	"f�$��#��C�;�(��W�Dq�D����^ت	�b�bzc��y#yE{	��:��ͣw��o�po_V��9�e7��@$4�R��&�[�),�S��-�+?�فa�%`��D�u�ϥ���B�s&�h�pu���Rp�^ǋ+|H�������j=�#��G �o��C�+�F}4)}�刘�|�/�@=,]y>��jg�_�A(B��������
-37�n�..�j�y"�#g���3Wq���>EE'�nA1.wә_f]-���K�%�C��	c;J>�H�TA3k��x�N�o����kT�n��8ч��
�^�X�֛_�.��%�]��F&�Ui����*6.�+?u�ȣ-Z������벋]��DH(�H��� �@�����ݮ��Eݟ��U��,��O�	w"nv�I^R�v�>�ȷ;=&g��(H|w�� ��9$z^���������_\��Q�y�X�4[bp/X!L�PFږA�Gw������u�ϛ��� �[D ��`�:��i�Ar�0>]�y�x
�q�B{F�	����ӈxS�Z��:���#r�l[ܜ3�3e�����i�����g	���[C�(vq$��A�	7�dj	���E!���t���4��p��h�|�F�j��1�F�+��C
�3�����s��2���}q�b������״,���.0����W�ϝ��L�� �����`��
N�}@��&�I������_�������@���0�B*�S�4	� ��"�9�/Uϙš����i�f�U5�֙Ď �*-��R:%R�5��t9y�*K�	�kś� ����~l���n�7��X4
�*�Ą8B�}�8M����ږf��e�o���X��2 c2)��	E+&��Q���Y�_2���0�o0�V|��kVn��)ʽ}����Ƽ�DT#�W�Փ�)^�r�瘹�����R��L��)� �����W�S'�7��X�`�Vm��V@�b�q���%���:�n��-*����2�Kx�R����WV�7�&�+X�_��8(�>�g@.��s����4#�Z��݈K�a��[�����OmCߐ��oN�%��Lt�f�A9����������	��h���9��QL���Ř�ǚ�=~�Eo)��]Z�����Q�d�399�����JX=|*݋� �{F��&���iY�;�pYf=X��a.}K]�}�D��-3.,N�&]g*��B�/���4��lQ=G�� ;�9�)�N�Ďَϳ�R�����q�����l
co����Y
l+�f"�8���J*cx��'b��w���x���!��P���(������.��C��C̍�=։
F4���	�II����������}#e���x�H��+��M-��e���:g>ѣ޳x	s�W�P�DNfm��X�:������Ҩ��݉��7_Ҝ�S>Ff�caZs��eN�Y�ܗdD���H$�t���X���:�R:R؀�?&8��L�Cz�n���ڽ&*�n�|�8�Z�O�Bs�8��i����,(n:�F%$Ђi�v���4�dk�wA��-Z���^S�����6z��F͉&n�i������x�Y����O�k�}𭸋Y;��_��r�z?�2�K�Թ�0�̏G�x��� �U�[��*��B$�Z�6'/�ݾ�cΡ�)����E���j���E���N��|G�?5���	.���.�d��|�E8�� � b��L�c���	��]U�z��������ρ�/ᅥCg�Ǉ�T�**��BG$��f��%�اs�'P��-G��?^�zfDC��� �m��Q�d�0�#�/���[ �H{���D�ҼSX�YoC�p�fa�m/�&^�����+aV���86ۤ=���cŝ=(@�3Rh��on:�TH��q����p�|�cX`B�0Ei^�u�\A�A�
�=�g�B�ݸ��2������7��"�Cl���C���t���\مݤ��Z��%:&�`��(/��b���Mz
P�YX�Կ���
��&����MY�mM&�J_����7��{�r��ؐ�&���]��n�sŲL�MH���0�"���v��u6~�)zm�,Yhb�E�Axh�K�V��Q�j*:v��^61=S�E{-��n�ݿ��-Hv|�v�+lQ��p�ք��@}��3BQ�,\�Z߸U�J&��;��XQT4R���2�]X	�޶����!:�hᝡ��'���m��Jh�t��-&[��P�Y��u�'�j���}�}�ł�jIG���)�o��p��X�[�/��l�c�G��rf)�I6�'�`�o�\���9g+�p��\���D��&L!�R�v�6�ЙPq??<�$F"���Aُ7Y�Bis���tYD��[څد9�e֏�Հd<�ky�"K�E];� �@��	"��v����S����A��ܩF��跳����ֈ*\�!*�'�GG�954m�9�3SMp��ŋ� O>�C#1�%�,mS���-+!;C���s\�4�I�O�,��D^�4�ADui�^����^��r����G&�9�0tqhJ4>�˿��<~u埗�"fPZ9avW��h�����p�v�#z���F�w���ڶ��Aħ�Y�,é����"h�̼1� �_v������ԌFN
$�{y�H��s]򬴆}"ڸ��i7��-0�x���\��bR`~�=�H����ty�X��H���h�6)��<�%hN�(���6|e��n�ĉK�a����rUFK��p�����9��7A���d���XTRX�3;A�,4E��w�����{ˆAx.`n�6����7��:�F�g�'�X�Ne����2��
?�?nY����()&Q�����7�7��,C��P*PW���q'�+4rPR��?�����5�h@ՙs�X��,�6��kh�3$y�������J�Xو&l#�=�W��a�(n���.��8c����3:�Oۥ#�7��eO��f����ax�;6�����z|��{͵,��ʒ�L�>?����E�T��t�@$|�D<{A�x����F!����A���*�c�ͪ����iW���:\���OO�(/t��ß�?���(�9�n&s��P���J����9~Y�X�>ϙA�T���P\���B׾9T;���ݍ�G1	'|*�J�@<c�}]�0��w��j7�«��QED���W|Α[v��O��Өs�iI i}�?>��<�\֫���?sf����u����K��%,�m�����>�p ��.rd+�~s��HR6�~l'I`SF���5SdJ<^�v���$߫�E�Z�DK]>�u�9O�/u�oC�-�6�jS���G�olJ�#��QY����ڬ��@�r��^Ox>{ULy�x	몏����G�q�֭�_��@m
v�m�6y�����^Dt'�b-��"�6P��е��OqbH�C�f���[3�UM�xJMD����j�+-jH�D���V9� :�Vk� ���v��5	���H@�0a�*�E����9R���p��#r�x����Hj�٘k�b�I�	j���1��:X1}����::1G��'��"DA<|�A���˃$�V߀�4e�\��_��w�.��u��,���S>b�M6[�6K��<��ϵ�ô8���!(��|d�$/���3��_P��A�*������C���ϻ�O8�~���8��<էCb0�A+<v�T$��0������z=wH`���3u�&�a�>�M�~V�s����5\��u�ç��{�!��w�j)���+4�' �"uM��6k���r����D�������-š?���{�{t��
���cap���!:o���G�[ZJPA�Sۨ���JĹ��bA����E����ؓH�e�X�:iڎ��aÖJ�of��9�MmU=�����_�1@�nć ��^�m� :~J�q���YGa��-�{G�   W���|�5)*l�G���W���ff���10�jQ*����BY�e��}��*�8B�䗬��8�6��v���/ۮcʤ�M1$�A����27W���$�m���zAC!8 ⿉�_U�t뮖���v�	�,r��h��ַ���DF��;��ǉ���Gb��ȶ���U� ��$/:Gk���te
�_GR4q�X���f��� ?�s֡!1��0k|��cJ> C4���Vx��#�kȭ�
Q���r��k��"��IRoU�����=i�r���P�Pk��eu>�y��j
/Y.?l?��ԯ��[:k��_��i��
�뢮۷N�����'��,^�_�t �0�gl[EH���,.ۂ߃9�9��7oNyI�;3�X\�����ki!�o�A�B�9o��o��*��:�c)�۹VC"�����R"ETxHfA��J�;��n��z��W�){ۊ[c��yV���UѮ��,[�B	�탵�=7�/תθ�.O1<�ɹj�	Q��!j܋��u�Nk�7tK�+�����I��Wj=@�x�GRh���2(/%�X{ek��C�<v���ui�)���t��_α�N�IU��?a�
�y3�42���?4+�_|�#������a����j��IG��_�`{�6�MZ:aX.�1̆fV^��V�OA~�.��4��V%���?�&�5�&f���F�x����_��}'�ӺNEGKf*7�h*��-��c� e4�ci���j�9���`�ED�֏�G�J�i�pdb.S64��Cen��iQ�B��T��tx��~��z�Vf���X�L��C�Tb�H�M+�9V1Qt �S�q�F��˗�Ibԍ	��(u�f�b��5�6*_���%�z7 ��K|�[;�D�V���H�?�{�=�$~Yuq�B=��7��4J�*V��J)x���Gpj�k��s��TG5(�Qd���+8Z�y�9ץ�Q���V��c�c�1����FB���W彁e:���58��~��?vV��l�1鋓e��9G7����	_@B��мKt�+N�4��$>+��AA��5���y��W�[K�q�E+m.WF���W�B瘍K����n�:�c�ܯ<<���2���r������=�;�8�.=�������m1�\_ۜp Uˈ�mp;����5E��0��#h,W�;e]����6L��b��P�HK[:�0C>�j��s��6u��i�#a�&�~�{�Ɓ�	"�b���v՘A7nO�M�C_��"MhFiZ��G������W�ч�?�#�8}O(��
r���T�DҼ��F����5xG�5O����
��Kւ1���ϳ���
4H]��~���ęeN)�׆��!Bv.+tzK�^�[T�Jw�7+���B���O;�'T?�7ՔQ"��΃��ɐ����"�C���Ǯ���B���!H��m��K)d�s�L��}�� }�G�ݿ�E
)O�ca:�J�2�ۥXn�)�M{~��f�7��4!�e�����@�z��4Q�b)��4�N��c��E���>EW�?�������E�5��^-��&���(Z�2p8Ù���O���]��N#ė���ٴ���\]x��h�"�iq�)ycL��{�;���l�����S�;�Q�����:�-Q��O�u3w�U�39��o�jP6EH_|H�֤\5����xŐ*�_3���6����.�O����TԎ`.jk�V�%Q���kxL��=���8�f�g��|��1��Ok��\��n.+xǏ�TA+*j{ki�ɴr(L����k�$��c��Zt�2K�:��#,v�@a���S�UF���@�~��HE*��x�T��;�g��?�],�i�^*$��TY�;�Ӝvby	?�s>�8I'��x$�Z�ͽ?�:�a?�V�\�u�J+��Y�F\�t��e��^1kb�O�=�m��"��ɔ�J]�tPԎ�`lԳ�/�Q����-�+46�u�J@ �����C��-��X�O�fk����+�����%%@~���ȳ�����BL	{<̤R�h�8��v�V�ɫI��E�@���I���@�p;}��N~�|��
F��Ӡ��Dp�:�U%n�Q��FѰU\�!�vnB=yeV��~X<욌�H��q�-�L5[#l�9*%P�ё�ᒼ2u�#��
�S9(���%w�����?'p�.J^	-#��*I��nW�h��ϩ�����}.�n���n�R}mq��$�.x��	͸�^�k2(��|�T�z����������_��~�Z��y��S�Ȓ<��{L㺝� *�5[�}R0���xj����B6wh��mI��;i���[�lT��d�?2
U���P��Ĺ�))��H��(S88�_D��aB�b���䕕�$l�!|��uO��6%@B�M����X�=w|�3�	���޿y�A�+�Z<��E�+���=ǩNO�r���x�2�]c��,����'x�0�J�Κ�G��.hs���*�\���?a�t7��������(�7���X(m��QC�le]�x����i��!qc�b�g5#�������W��=����u 1������eO���wu��d���b�C����ќ�δ�~��r�b#d�v	�|��6���Qv��[u[5������~��*���(؆�~�6֑�Ꙫ�ꑰ��@���](O�Ϩw���!�����G,��3d�����λ��/��W�J�I�~m��Rp�:����fY�cbv<VS����v�]Β���0�fzƶ 24���0��Q�Ca#�ub��#�󪹑gcQ�Ő��/s1Pv@��f�g�*���-j�T�@����{��k�������M��������6R��S;$?�v���a�S��H�aK�2����7د�h�U����R�S�2��p#�@��P��_�b���b|�j܇C^�kր���)
s��\�c�3Mn��.�U͟vl1?�y�Q@ yoK��� $�P�V�?N���Z�n����o�hjz�56���}�?�k�Om��o�K��e���;ߡb�t��lj��U�?�ֺx_�}��G��r��c�P�d,��P�e�W���`����8C��������hS��{��[d�����A(�ܙ��&���cЅ``�	����9
�9������Zշ��}EUi�-��Jε0�xJq�&���"�=�����'�<��z��{ �J¬��	���T��Y�5q}*)Cx��T�3�u�ރ��V���TW�D?��(�z��W|��( .Ջ�$+��P޴j�,����f�1�@}��߂=�	]>Kq����H�Ē������H��/K��,�^Y��O:�)���cJ��/�BaVƺ�s�E^o&V
�9�1R���:{uH�>��rߢ 6�<M+�j*l��N�C+����h��+�C�Y5�$()6#�FQ��7��G�c��UŮLȟ֌�ڬE�s,�W��T9BN����,
��Z��/K0E�%��#�u�JU��Ty�PYe�D?3��5�%@�O;SB��kl�z4"�l/��A�0|/ra�xk�{����e��F_�~)7��Q.�~c)��ǜb�&���*\]u4*rS����w��$?�0�V��O��,�k��r����)��WV�\w�NpKT]��J�h�A�}8Xp��uw��ͯ ��������8����/�rR�
�R���4;oD�~O�.&�e�B&���Tlw��ο�����$���0Th/�x�/�/�S�Ƕ�z�H'/>c�Z{T�W�&��?bܯ��t�WO�Y�����ߙ��b�L�^w*���ϓ�V�����U���*1Mj�3���i<!uf�o4�}�\��c���ZCa�r������=�wp;(컙;�����uN�nN�~M��16@�t
��	� Yʨy:EBۇ�k�S�j���vU�Gع}��'�.��VU����7[?��>~x�B��'�Zj׈G讼�������T�{[Ρ�\/�ɤa� k�o���m-�@�� ^yS�����-�
���B�۴���랻$)��П~$vR6	
��m�DWM!c�q�|x��Ple���:7��+-�(!r*K��<����4+hR0*!���=z�o�dL7f��J���Wv�&HC.I����`J���cW�Ph���x�X���+斜+@�FBf��Vv�X����l2����.ۧ!���i�Kz�J���|?�Ѝ�KL���vI�Nz'��]P��>t��Y��)w���TO��E㜃`���]La��|�6���P2�|a�B[�,B�lJ��������no~�ɯ�����V� �6��𢵆� ��=�y�n\�cPM�V���j�@����we���cx�
V0~�c�f�~�n��Zg�`Navu�T'�-)`J���軠��4DY���|.�R��y�(�n�9�Ȕ3h�d�F����u-�)4E�>Vy�v|��CZ�Z�Q(��Vң�:	�a�#{,��q��O�P�A��ԇ�<��	�����d���r،��ȁ�����UI~א����$��~��X^8:}�^,?����c����AƑK�dg�7�S����)0.�������@����2w��H+*p���������X꘻ֈX�o��V�O�m�<�T�,6�D�0�N��eS�ݷ��M��ʧNiy� �j�$��G)J�J��O��k�2�Қ��Ǎ\��N.+ᣆ�?��.�f�d��f�?�#��j5&?mh�avx��Ԥ�-b�,�3�m ���۲�O�b!�_b̴I���{��Õ@=�4!_�1!��b�!��ŧw��A�߳������I.cz�&(���D�M�����@��@��b�c���@�Mxp��2jT�qm����4�J6,}N��X�/U���N��9���,�t��)�����n �}O�!p����^%"`N"tME�wj�m@�e(�}�m
���g���4�C;{�
�������[_ ���JHR��u��*��A�T3,��Ļ8(zP��U�A���۟a�pO����ײ@ ><&�Í7Qv��D�"-
Y�0}�XKunY����H��͌e��z��ZOA����a��gt;� �(�4���eX���|�u~>�;�%���`.�,{��N�0���均�<Q]N���禑*�ͽ�n�E=	-���zN�#��� `��_e�uw� �.��fn[A����-�H`�8��iw���gmג����~UW�����a����R�m=y/V�	���[�m����,����w �����k�BU��s�gӰ!3�^Q��G�n�0����'�r��S9/�뗪�и=��MXK#�n��+~;D��`
���}����}U�/���R����cBa�����HU�^1�� �Oʏ�[V/��`����_'��R�NW[E[�O&�êf������Ϩ�2b��1��*KF��7{zJӻa�r�U����z/������b	Bgˡ�~1������wy�Qնg��5;�*���c��58��T��k\X�~c�i�ɴqm؄X�hD�v�X6�޲h����4� wX$X*4�(�B�Mg�{���y��5<'���kp$���I7�����<��).��[>A��:��0�`��y�O�iX��n�m��c��:�t.�s�+�vtCA�d��Ђ��R�괂&˿q��ck�\ 3=�7dum��Qp�R$���������`�T�/q�>g���U���C(��6�~�3Nlk�����7ٟ:�Ke�t��L{���q�W����`-YMPp�v�	j�$܊�2�*g3�o.���6��jUq�F�*c��-�V�c��K�a�i�C��(A��a"�\���d�Ѷ3\�>�����5 ��U4��R�����|y�S?@1s�.����C�6o���*ܛ�.��{Dg��j��3����6�k)�=c��w2�6b�a�ڌ[�G�]͸Uխ��wa#��X��m:P�@wG6,'կ����p��#5�}J]\�`Io���	�|�Sd�
A�d��H����\ٿ�dkG�ݮ�@g��\x����n��UZc�g�6+��J	����s�����끾�rr@�LowW}�EI�YX��8¡x�:�p±2*@�N����ʻbP�a��j���*)G8�ǲ�E�A�'��Z5�f��ӟ�ZC�(݂�kơ���s)�W!�� &E�54,���?C�}]��w]]q�LT�C8��8�/BA��Yʽ��}�����S�?Y\�b0B=�p����D��H5�������Juue�I��m����=q��Tu<���{r!��{���n�������#9�c�v����5�XrᨚP�YĢ�U�{9�%�I��������W��_+�g�����:[�BW�C�1q��+7�~h@�^���Ê��Z��:6��?׵�5��1���O�x�)�MCl�K^%^�@���xWV��b��6`Ԗ8T�I�����'�ȭ�����j���V_�ٓYgV��iq�e`�ɿ0�ql7*���Q^�axW!�$9�������RY�qX�WV�8{B�<�UC��m��7�[�P�y$��$�:���S�ϙ{;����\\��P�Ut���s�e!L�J-��p�a�ʜ�[
i1�0왮�rm����GvU"�_��5���+���H�y?��U�8�b��`vA��;����lt렓�uG�<�af���Nn@�2�0��ٶ,���G_��J��;����8��_��K��rN���70�F�6�����[2Qgy3*��G�P�a��F(�x�ޯ#� f���=W�~��P�g%_Jҡ7��n7��%s�P��3��j�T&��"0�_�
Afo#�92R;��^NhI��?0K�2h2�Ev�o=n���"�t���7J�0k1�tf�I.2�����\�Ǚ� s�_3�i��B�r���V����i�1>s��XV0 1k�)8�bE�CV��E�=T�W��O��>h ������l�C$�z�b�V+�BRx��p)R&��5n}��N��W��~RR>n���}�Y&�.����-' +@\�gS6,�
e��d��T+�X��M�&���K�9����Wِ&��K>�؊��N6W$�ڼg;��MA�/k��o3�����!L�`*���v|�6W���Y��u��-\O�Zh6;4gsR��dA��'��h��������D��HsɃ)�Ҭ��u�R�&���K����R"<oJ�U.w�Q�Ǩ�?�i����,H!r��K���?b���q p�����V���]��n8�#���E]!٦XS�C�w�'~Ɩ�7t�f��
�v\��x���IMlx�5��$�9����ew&�cѤJө�@4�K��zi�� �fX�43u��DM�(�\�_ mK����|��&����)�nٝ��?�b�濉F������w�����I�P���Ly8�FlP���-�T��� �(���� ���D���`�����c�D^8�֌�_�:i�)��.<�Z��`��C'�3ͼ�]��=��ӗ�dYMs�����/gj���K,� I�oݽ�U���W�%�\�}}�"�OQ���Ԑ�c�E�V��F��DV=�[u�s��_Ǆ���������j����z9��Hd�{��*3���e�)_�R:Op��h%#R�7Ӿ�R�[v���1�����`��6���#}����a�֘��y�@�{��%'�O����E�͕R�j���NP�Zf#N���O�z1��cD��^7�U�fD�AóB�E�F�i�2��:`]~O�]ǿ���mƈ��E$@U��~�)��:�F=��'?
)�������=� ýa�� /�A�E��֞������A����z;s�y�3t`M��cUkK$?�\���`�3�Bu����E#��x*f�n���zhV��m~�C��\i��D�Zl�����bu	������G����?��f��i�Y��<�Q�gy��ص�*^b��~�����*�>f�2;8B�T���Ri�ߙe@�Jg�4���0�-r���%<@���Ѹ���� �f27��r����{���le�G���~f	�ï�*���u���V�_lKHJ��6ʘ��c��=��a�HAUw4��H>m<��GLI���d��ru%�0ቭp�JE�\��-dB<�^�F��gj�a�`��bC�Yj�%�A`=������b��C�bw 3hE��
�g�<r*utu�g��=@B�W)�Q����c�E�=fY�gKۮڦ��n��J��6���~��
kQ3M�ex��ãP���~Ly��ȳm��@(c�e<��}��D��nu@Ը�>D��� �R���W9ޕ&�K�:���W>>�8�Yo
x��z*�:p�.���a�_	:�Ȉ����:�	N�?E�����n}�I���Ϗ��Jw��,�smƁQx�E���^��@◴��:ۆ�$��\��a�Z~����zap�o��L�������Y��VVޫ}\q�ǪcӘw����{�����ߎ�D-f��%��7���kC��׷:Y>\{^�a��J��.&p&����:��}vK(i��k��`�����oX��m�w��@�c�47M�B�}�K�fĵ����|W�/�W�rt��I���h�UtH@`��OJ�:���1k�r�D/��]�80�Ac��rJ#��f&�`�b��vVf}y��w�XM����\��D�kå������.��ͻ�x_�%��a&�t�������G�+Gl��7ٜ�̵��}{n��sZj����ؗj�'�#���+2����}�s���r�p�[B�מc0����뛸��Y�����s�{�^�����{��U�:	`��Lt��p�8]�]�������:�S[c���S�y�� )T��;6RnF~ E���R⃠Y�#GF�p>���j���A*���Ԋ�y+��$�����l��o5���s�<�#��٩b}�1(b�V��+SC;և)�$(�F�M��?�<꼰[&��k�h���Q�!���*ؙ����e���9ʨ�p�36l�zfD��"��ba(S���.K�^>^�2IM�V�ξ��/\u�$��Gb����3/�5l+G��ꁭ�ͳS�e<�_����>Bm��2�n=�1���e5�@yN�R������-�e]��e��8jp���G'�~bf��LHl�<�i�9a.;+r/�Wn_�Ki�ʍ|�|n����[�`S�YT��к[�b��J��D�����m��]�?������?h����Q����m���h����L��&��~��k����?�vP���:�~��Q)����bV�$,,��җ |�C�K�t"Z���46#����OHDC�\��9T�-��P�(�:�ڋ�㘚�ι��^��>l��:b�@b��)���������[��z�6��ǒF�kWŐ�E+�o&�:�fjR���{g5��`{{b]0��T�x�'���AG:X$k�x�~�6�q�<��q]�4I�,��D��C�䮣��R��H����ye
u$�.���ю9YI�P��*TSG�eE�戮f�~���'�H��A����Y�9�5H^ǿ����˞�-�M�#���Le
g)3/G�}I�8���'��}�g�Nz��k,�YVHњ�;C�u \�q�2Rʁ�^��t���5�� ������է����3�D�S׶㝸ś[a�V����J#��4-h$�Û��D/c�b%7=T0�̘Z#p`+��4�_�8'�{s�Gn�{Z�|�y��'.��:X{D���=(�Ɣ6�1�Fda�9��nR���·�7啐�a-C���!ɷ�G�XU�����)}��x�z>���|l��f��Uj+_��6{X9�N���]�I�G�"s��*,ZMe0�9RA���ܑ�2ozEp��|WF2?Qϛ.�VV������eX{����`Ћ��]\ֿ����]��ªd�F1xB���8��0$b�/pPگ�+X�o=������}���pk��j_cl�Ѹ�>º7W0��,t/T�M;��>����9�I�-�Н�,j��Ù��D�@��[1�_�Ct?<<������������`��9��9�����+�$#l�H�H���W)��&���K��cq��`���"�#��Dz}���msE@0f��(��`fW�t��B۸$��nO�wqQz;Q�Ѿ��{x������x��vh�G�/�knJo`R[��F������Y�p�w��+�2"�Kq&n�먾�lU���l8AӃ�*XBvp�>�Ro6�}�~}J����:�y�@�Eq��֑�C|<�LG���+B�-v� #m��|��s�1{��z��2Wh&-ߨ��2�-+Q����CĮn�Zn9^6C~6@�g�E�`�ͫ��`��G�E�?��Bc�{������Ye~?W务`V� ����;����v�&�Ej�E��-�um肙RROK���=�ɟ���;xx�6eמ�p�ElyI����\h�a AK��S�|~�buQ���j��꟯/»�j@Έ�s�����c��72{���-����D9�Np�6�M�����qQ4���	2��rL��R�{
w����n�h���|���G�إ]�`l�����r�(�;�]�m=׃ag
�"��A�NG�E��b�"�b�'�syÄ��B�C�G��:+C�%�f�i�^��ۗ��4p�,8���wh�}Q�|��>�#X~��-�h�XPx��7z����Dd��F]��@��ш0(Tw:Q�_�Ȟb�)�R�6F��Tc�ߙ9�q��=�\�+��FFy�w!� �L��`c��Ĳ�>cf�9WK,i�@�p���j@��HN _xUc4kad���?VQha�AF��J@j��o�iOb>R�7U�*�pΚ��X�:�w��$\�X�J)2��nt�E����傿i����T�<ʝZB�HUd�0yK��s��v-D�W93^��P�bN��D���G�M|Ν�A�?�b���3�ը�w�s�n�+��^n�
!�d�8o���7H D,��Z;r��ӣÊ�Z}?��6�\�j�w���g`Z��/�v�ih�`��.㬍3���>h�"��,hV�Lhj7�� �Y>������c;�A��cVv��^Vp�R�d��A�^B|.乶����"�O�<���G�����߃��hFC��@��bC�O�ꖱ-Uk5B�z�Fo�Ǫ����'��E'O�_��8��M�rls�8�����E-�t:�.���\T�Q�r�i�50�W��1Q����P�q��g�r:�{�S�,U#��6#4���.!��FT��r�BJ7��� ^�M��-����R��X�ILp��T.a5n"�;C��rg�t�\��X:Ae7Y� H���6U�}+$7T"3I�eΗ_��^�7$ȧ0Wc���E�xo��l���Ms�|h^�6�w�j��6��%w�%4���ĸ�-�֤��G��������LE�k�)���P�SC�7�%��?�;JI��lq��ԡ*���A�vp�j{�~���K��3u=U�WC'f�����+��� ����(_��2e��=hY�M��p����*�� ,Go�2�(nl�����x2���"�}��v|�oPU��.�5��Ļ}���|/jݡ���i�wVV%���<�}�;����?B���}�0�PL��ԣ��t/%��8ޡj��2��n���h�0�-�&��_�	^������y`Q����a�u�����9H�hY=C�?��o�I!�Q�DU�>g&]=���À�$k�W����jA�x�����r �( �H�IVߪ���$L'��|�@RZ�f�����9k����J˜���SL���;G:^�����:6��5��ӂ4u�5��X���1F'���RM*�I��:{k;����\��{��{Ǹ��ܐ��L\	�Uu�;�X%�c��>�����'X��m�L\Z}t��6�vБ�X?�nš��+�|�n�D�&4EࣂI>�)���{�&�p��*�d�D��G��M��ph��x2��5�P_.A�>���~̩8Ns0�� �߰Yo"_~���c��)�R������"�qn:8��R���0#B	��k��ɺS��5�'��w#8?�U5��8�M
7U�2+�E�����8�\�-^}��0|u�"�N)&,���B��o�䡼�J�/��:�%�5�|ː7�XU6b�f<ߒS>�%�k#�:ٸZ�N��NI�O}`r�m^��X�D�M���Jx� K���;K�F��r�a�Ih'���}G��~�m���gƘ�c8 ���*g��J.�ʍ�{��A~����P�|�<� Zr)0HiC�5M�/�9t|� �3�cu�7 s�h�e)zԞ�E���&�u��X�;S�D?�v��KĒ�����h�������y�.򿿳3;*�@�y�|[�3~�$<�1�KS�g����1��D^	5�1{H4h���?����%9�ԍ<������<��^;~,�1�=~�#��=u/�?xS�M��Y���+|H����u��E�"�zط��@�))X�K/�xr�,ch�����j��r�G��*"��T�Rp�z<�}STyG`tp��MV�E�W5TE�iۧ��������tx�Cظ̻U���#�����]k�T���k�l$��G�8p݊~�A��	Z�vO|������VW.a� W��1��AK���̰�&���9W�6�KBΨ7z�N�w���Z�/�( ��ڱ�Y<9#�*p6��6�nt2A�t�4�Q��LN��Y�M-k�ՌH
����]?s�,�k��qy��!���١�\��g� FWH1c#1]Y�y�Z������;+�'`:�I�qI;�>��L=��;�@8��xǟݹK�и�����]�Ś���\
��q;4C:���M1�c(D�c�J��C��l̵L��~��v���cmP^�m���]��#,�z&��U�⭆�p�C �&ͫvK�;ɦ�`��kɘ�J0�(3|i`7�"���vqTb8���YǗC&\Yg��W��A@�����fs3�!S�'���r������l�=��ty��>t��;�B�zO���j�����xP�˩���
�`���XuT��7zG����)��^}�����»FA�j |7�&�ﾄg���4��A¶M4��S	���u���*Z�c�̓��OE�׶�h39-�/�ȍ�.�T=�/�F=^�W����R5�����1��R��~b�� J� �U����N�ttS�G�z��l���뎱�E����::�'2�����M~ydN�.q�tHGm�v>GJ�?BoXU�l�|��2�j�q���[��߁�����X�w��d���V��;��#���>ڿ���1P��p��C8�D���֐Ed= �Sw8Pn�}A����Huȋ�u�֩��Jϕ���o�r��<��%?��	� ��0�,<�����#N�xH��K�f�ѽ��������*�G�÷57�N��X7<�.��PZ��k?(�hF����b�P�<���.op���ò�Ӹ��L�
F�W��R�:L���!W;��v��]����a ߸ ���6�;З�r�coZ�ᝨ��,e[�;���ˋ<���ǐL�C�u��2z���n����X�7lb�0}����+���Q�0:N&0��A�V�����l����o��?aD)�贐'
�&�A����M�R>K]} }<x�Wg'�v/Q�Ҵ�.>��ز�E�<����K^�nR��R�������G��6tլi���@j�k�͸���ь�P�s�`��r�m�k%4��d��=���t	6�-��~�\x�_�蟦�Qq����W�$�o�Ba�?Q�5���qo!(����Pm⣽����){܃s�r¿.���bY9�(<�eE�4���Wq�h�ܙv�ú���o"3f�k����Lxǂ�x�Q����^B�o1��[��v���E�i�����$��SE��
_�f���3Aᔚ~B��n��d�mD����1���[6�����"KDHl�;���V�S�|�p��{VJ��=����L�k #r���t�
����go�c�r�<S�7�S�]�rL9���� � "T����jH��D�'�,U�7\�ȹ�G=�-Z�dn�,�I���]*Z,N�㩏�iXЀ�uƶ�h�H���5�i$_^��t�V� l�h�(H��im/������Cnc�Fh]`k%*&�G�;n��t����n�(i��$�?Ƈ<�*����Hn���7�u ���:��RAD���c�U;�f%�I��	R[$?�W�cr�hڧ�]�N�$
�.1?Yy��{8`��������쑊N��B��E���k�7$p��*��װIT�槛|:&��C�n���@)V!��{e^�H��'>߶Yv��9Is��P���cӨ�t6��C�p߽���rGHw�l��b�b��������zc�oXm�+@(�	6��f�� �#��j����n�.�R�D�K�B$2�(Uw�D���O�P�p"M�U�f�^���;�}?��) h������Xj��P갅N�D�b�&�F<O>�ss-�+Y�/P�,�q~u�/�j|��������d��a���S�n�cxr<��k��\��l�OLl
���=cY��=0�O��@�\�)�l����.�Lk�KH�0�r4SAqp^h�P�ȍS�d$�n&�ԏz?�>a-�lt%K���;�q3JLP�?n���3h�#x�ƾ:Ŏ�H��zgSF���BbY��P#���+R�_���?���}�t�7���&:�p:[���j����G�V�r�6݀50C�������7�ՉT�6O��pz2�h![u46fu�0Җ4[l�K�<�7AZk�n���q�7:�^�T��»�N��+�s
;a\�����ܚagc�	Í�a@}�5%�r^��~kd_{�\���@θ*�����J+�F�[^)����L�k�K�I�_��pj�İ�j�n)M�!���H�s��AX.pDF��
��;���IcSL��u�I�."���`{�������-Qy�y�g�؂�1�@{r�xvq'�H��4IN+�ۼ�_�hc��nox�c��f�^������A�q^�?M`1f�4�����K�<0�4g����K@t��LV��vBȟ�魀�ð���[�3]�?~�v\��4�0�$��W'��y�,HM�e���`�N�D���4��1u7h�b�;_�J.�����K�5�������������/u�]6��Xh��α�ihw��L@�g:FQw�er�`̖��#����ѵ���:yC��:�Y�u^}y�87Y_)�h#D�J��جI
ړ��1͍�bz#?(Nbsy�e��-d����ѣx��'��kH�4K:AXW�J5`=l�T�O����w�]@�"���r"q�H�k��p���q�V�����\ܯm-3�O��T40Č��œ~�aGH�fk7MO�8Ӷ��]N�@�Y4�hx1���Ś��9.����3�^��=-��iNƇ]g꿎��\'��ލ7�f+�8`�"r�Li�rG;�ӔC�ZA���}V��6�@�9�a$����[���kqk�1P�����"ڗ��%��{�]^s�
�25Z�IX�'PC��x�q�j�t���� �u'A:)����٘+������˚~G�Sĥ�ؽ"�
��N:��<���zP�r[��Ui�n���G�f���x��}|�l�2�@���:R�0+�%��nP� �;� �׊2U�}�W�Q��$.u'-e�sVob�4�"�:�B�x�t�%Z��y4���$�O���
X;qe�P<���@!��b\�`���<�-F�A�y��'�v)rt�'�jF���o؞�J�	"�`E��"dyШ��5!rP�U�"К\$x̧�۪c�yħ��p�IDV)9.���N���b�'�Ԙ\wPj�d��Ɗi*�JD�},��o[Sٍt���`�I��\���D���M��bi*��·z��d}ŏ��f,��1?�8��ݒ���w`�ғ0*��w�"޷�g�k2�j��ʳ�|"H:���K끼񱲸��������)t��y��Vi��7o "pE�������{��}	�q���X#D/<��.�{��\�_($κr�j��=G��/(u�p4]	���hM�I�S?�B�Ed��Wt�F·M��{��h�l�L��"_W��*�%�0��y��� �ur=q�>;:4f惞�!�^e˅��BU�8ܙ33�j������whC:+},�mXh�
W�u�t��H���&����?O�!C4���湿�	ƛ��x��ᗲ�����-x?L�lm5�8O
�he�����+��m~�&��yRk�߯v�R]� Z~B.�3s�H��\jG�j�Sƌb_m3,-Y%/�!&�qv�:l��$��$7Ǣ��G\V����_��~����ע3�C���?� q��0xc�Cqeg�����{��D�C�'ۨ�T�I*��p����H��)��w�Q�Ţi���j�91��Dfc��K�t���o衕����ﰳ;c�����t�Z,��T��b�$"W$��`,
�<����G�;]���j�v;ޓ�Ĵ������(��ۦ;������l3!mK�8)�Ѝ�9���FJ���h����s���o�(:��B�Q=p8Ӕă�Y�''uD�/���I(d��o�r��"�KA˺�f�[>�>�EJ�P���U�<q�ڊ:(J��H/�(�Hm�8�'����Pz�
�)�'���Z��~����Eh/��~=��ayqriz��,�]A _����5@]�oK��z� ��>���{�� ��k��D��V?�V)��1Dr�� ��}f!�kz����_�5�c���H����4]N�f�5�#�F�*�y����q kI˓W �P�SJ��~1�bz�}S��m4S�i�H��rd�w���
1�IN�zƎS'W�T��:R��^�h���v�q.ɫ��\��<}8Wɣ["n��.�>�!G�iW.�4|�~j�m���fA|O\��x���/�ډ�r�p���{���Lc��tb�� ���=,d������xC�c�fBpڼ�^��.�%�ꍰ�~��#�F:"�UJJ����������N�m8������dR��IK��ϟ+d����tg ��S�&�x���){'� �O����E	��)'��[��?&HF�^�k�����9��u�oR�G�V1�<��bY��-lˀ�$lk1�ۧ{�P��Q���0}Ϲ�55dȣ�j�Npp��Ǖ���-��w��ov��i�b�pHM�����T�ڇF]O.g�"@?v����N:���CI*������Y1/�����D�ˮZ�\��	G같���$� =�YJu�Ev��֣�1�=�,�[�}�.7�8)	����$��W �><�I����=�^�_���Wϭe�pT��@���G�h��i#q�Y��p��.��,P����!����)�ŵQ�<�o�=�����k���M�mɪ��-=+!H�=5�Ӽe�|��Q�ϱĹ|:���D�e�0���\{�aq��0����`�&>,?A��܅aۦ�2<���P�lcH�l�l47�� w��E�]By�a*�T�n��猛�-U���"bV��0�7�eׂ��L}�&݉No�/���!�\Nӥx&�=��|Xmt[�r�V���'�Uo�q5V���r���Qk��M��D#ÊdXq������=�f�X"Qޙ�Lz�.�X����!hY�d��:1I���r�yg�L��!fW��+��=9�u��E���[}����nFeJZv/���1��Wn(�쓽na�`xh� KK��2zq�	 �l5��˵B�Ut�?�y�"/����8��ynj��%o���>��S��7XG�̝����tMsBa��N�D� �J�őe'���4�v��ci����R	cTǢ�T�~���ݬf.�d�H��v��2R-y�'�S���X�!�d1��Y-v�"6����n��	;�Ȓ�;��g��+����߫,��H K ��Vm���n�a7�<ft�,q3Ҫ��ZI��`�K'JD�2�����市���C�;	��I˞�Դx�E�b4�d�Y�~։V���G>O��4�S>FϖM��� �L�:%<Q��6a�� � ����%H+�(I����R]����}���\!�A�PF`��#���re�̴{kz�9�ؑ�޷�6��<{c�8_��影�EH�pT�`���,|��6@��~2�����RG�Ɖ�|����pf�f���q��f$�?@�Ca�!o~�;�̒��mp�ղ���=�I���W}m���H�$��t�����Ҵ27F����4��Y���y)�|���5h�7	'�h��#�.��u
,J�X�]\��y̲��o�N��Ů���Et����͟�q� �<��4]�1ş]�k�b������N������A�6a�a����c�|��1���纑D�uS�fo�uk�����n�&\�#���Ub �.����`��ü)�:_Ī�z7�zB�%�D�jv��:gmVQS���"�a��l��D��B��D�j"�faXe�\D����K3���u��w]h�E�i��X�!bJ~F5����CT|��w��̛D����.Df'�+	�����@������/���\��A���V��J��I�F<p��}\�l/b���#��ؙH ��]n�c�M����t	����w�L�9j�m��:G|���xrL c�.��I��m/L�"V3n(�7*������7��I�h��4K������Q��H&ͱ�������I�0�gf��2[��X}w�K;^�{�(I��Z9��0d�-��("��'�j���Է
��~*�%�:���1˽�S=𖖎��h���R��7��$��s����>�?V��U��|�[�5�n'���rJV�c�8C㎳�
|�n�L~V錮P&z�>����2%`B��m�!8�b�Rp��R�%:��K�{��e�ag�]��lC��e]Ts�ֲ��dL�������"	ޭ*i��V��;m��qB�Tą�e#��b�͗4.Lic_V�Um
z1���Z�߭eOMr��򹴊�em'h��e�g� ���GM�;�������@RC-X�DƠ�{�qa��ӳ�����x����˝�r��h�Y�Y�A�v�>K���霳��31ihR��MC�ĺ�9eh��#����Wi�
�K������UwnF���R���i���ˮ�	�L<d�ӫ���^�lXc��l}��=3�81�%�ȁ���0�}��-1�ô������+duk�-�=1Q$DN���s��?�������>:�8���JhIq��=vÀ��Q����1�/�8���U�q	w6��(�$��K�8��'�r�LX�z��y�R�Oy�=V�����3��@3�xau��0:^־p�N���00�.�3�+5u"L�k�g��'*w�Hb�'��i�.��b2Ob~��9������*ݯw!���a�7�v>�ܹ+����x��M�|B^��<j�m|?���ns�D�P��K�֚�Z�Fk���jJ��8���sA ���Fc��}��� ��g%���`0�{�5#'�A��I�o8$b��x�ڝ:��~�/j{Ag�lh�{-��81L�cO&��l]���K��	�,��.�-��c:s�&���7�,K\$��@O������՟Nu���I���4D5X/n6�8C�y��b�Z������\�4���}>�[��8;�y)�l{��>�bWvHY_�#��h�����8�!<�%�����n��cQ�Bh�d)a��/�*`s�ˌ.{��%	�Ouꕙ���Y���S��C��k�@�)��C�4:@6f�#A鐶f;�^T�B�x�$�N���b�{3�=�+^k�Џn�6�ob�>��w���c���Z�Y�i_��|��4��<Et�c�L��K��M�T|7doqTz0��Av궃X�WU�+�C-�����"��XZ��+O^`9,����;�-!lV}g�9
��!��o�}�җ��E�dl���-?źR<����Dy��Ӳ���9,�P��Fz��":��q�O��t�����Ǆ�P!�N�Up�\o%����e��d9�"��}��G6XLt7�+H��SMξ�V]!KYgvy�⅀�=خ ��e��*�������'LƷXA)'JSգ^��yӞ8�Q �H�#]��J��`�f����UO�-���^�9u���>#��Q�����gxB�%GS�l3"P|ޗ��VW��!S�^�mx�j��>�=0�f�O*R���O圭~S�{���/�3y��ƣ�k��zjG��S&��\�/�ĺ'W�.�_
9��@�w��U�3���U)�Ӄ�271���{�7U ��}�TrJm<gH��!�1�Μ��jmt�~�o��j�~!h�NA,SP�V��[ݕ�1��+R�$K\d��~�d<q
ɋ"JA-Z���b��m@a�6C���:�ݤ{���e1���������?>s�i�.��0��׹�U��.m��J#c"IU��J
�
b�25�D��c��
Z���z?��V��;�*ܻ���U�z�=e��0U�I��/�Պi�G�9ٟ^G!�,V�r�G}Z�e�N\Z�)�{(��Gab3���w�3��R�G�߰���:OVZE��
k��O�=��+��Y��>��i~�%�����ْP�׶��(_^�������e���
��U#�?�K��pg꺓��s��C
.��f^]��W��ᝑΪ��c�M��_�j�=E������0��QZq"%�:��Ğ�ؘ)��ԣ��Q�:T�TDȵDWu?*��͇��Ƭ=Jx�����L ������hB�_�'�SiԲ��5��	qKY�)���2_�m����z���dNנgW�F��\uV��L��ZvgJDSD������Z�����b-@�y6ji�����#;P���Y����H����.:���?f��4_=���������%u�"]Q�;�'7�wq�Lka9��*�}�2K��,9y����8��c����;�m��j��2�e��צ_D�D۪��+j��<+��mA��e<��4����۩��GSIV��Fp�F�S�$c[j
lV�#�h�� vV_a���������%X�.9Ѩ�v}Z����0��-�؈����Y�C�	j;y��0Ws�޸��� ���Xv�>̹F��_[`ڬ��5�T���u�Rf9���~>Õ��YgȘslDn;�@�!6q��@�yuԮ�;�
@}�#V
~�,w_id��5����y� =��ԋ9S;d<&��J�dKe؈6�$����A�kQ�� ��)}0r=Gs��V�����L�Ѥ���2;�Zlz���h[8h���(�R�
HX�aPC��W&�k�?�eܟ�-ě3�f���5�����FB@�4ԋ�A:��r:+��ޕ:8�\�Vy�ޗO]�L��< YG%!O��`��v�9oG������Y=��ԒU����gâ��f��ahM�rj4�(=��~ɲ�� �YH{.��,34���;�v£�SD��試�9�"ui�P�M�:Y���;��	�dN�7-��E[�/1��K�
a���R!Ui�V�!%���D
j�A�c}RT%8ȆyFu.��nYkП��I�
���y�oG?��C�sT�긽�vsdo&Vlp@%���6\(L]bY8�Ki����0p��dQ�e��n[��Lȣ�e�s�&>Eo��:������(�#�fN�s��߯���3��-��q����:P�����y!7ݬpi��&�/5��SE��R�6ie�f�n�B�� �ӿ(#�r�iL�����,���%jN�Up;�U�P~ڞ�m�I,�
�q�8��� �@���J�Uyj�T��?�D�c���L$�{�mB�v^�j�.��Kz�4�^��@�G}���X�y����ҒQ$�Tn�dس�+nE�+`���O@D1��x�g���|��a`p5��"Iѳ���[M�M�&�)���W�Bu�GZ)fY��1j_���T1<%< ��by��-80��aJ��R��>*P��aQ�_�h���6���K�)�x�c���s���j�Xi)�^�}���:Z.��)�������#%γ��ǤPi����]�����i�p���ҍלc%])��\��	w�qϦ���e�YDU�M��V�c�)"v>�� ���<.�o����m�ލ���G���=���qj ?
��mx)_�C t�)�e���s%R�fƯ�F.Ư�;�51x�@BQ=��hU�� �b%���$�W����6J�J+!��^E��S�u!�'{rE<Ϫ�1����lڶ~#v�T�44�pv~�u߻Թv�]���^����e�>�쭷�sG3���#쫠�@��\you5we��-#f�l�ߍ`�F�-��D���[-6a���1��U�4:�(G���ǻ_l���1ኩ]�����i��c_��}U[�1�jM�����H�-���_J֌'wQ*,7Y�[�,{%k	����>��jj�ļ����7�Һ�\�z�;Y��i��~��?Z�x<A�p2ҤF62!9���}�������݈�|OO��
ݪ_8�2@�y1Z��.D��odz�U�I�`1c��[<�ǧU�L*��)&b!3�N�� �B��s����2�S\2�!����@�V�7���\�[7�Y��"���z��M}���]/<�Ti�3�O���&]U��o�Ez������}T�~y�F=\��������e��>+Z��d �-S�|��������J��a�q��G��"7�ɂX�iI�\�hPC�ڽ�Y:��q�y�nê3���b�yO_���e�,Y��}o��&QD�&U{3F����#ɵ�1(/G�C�-h7�T�A���'m7[џ���<��[��`�L�4Qң�m����x	TSI-K8b��;f�x�,�u2����4�%�y=v���Ο�Ò~�!�2t��C���%���E�������h+T�VNX�'���He��ý��ax*���~Z�.۫&����3�v�2U
p����l&�������>�;������C*�¯D�s��!\|�	$�wU1|}V@�֣[h<�;JU��if6͏
��~Ja,i�7z~��W���#>���8������2�+�]�d�����@K�e��(���#�,�z���*��k�p$�L���_��i=��U/�
�^��ĥ ��Um���\���2�5�;�_��*W���^xAb2���?�W�>�r/�t�I�pܴV�瘶�� Ƈ���T?�3�6�4��B���7�pT=\�g�r1�d�3���f����A�wCu�Up6��A�����%�ӻ�Y��/K���R:�B�Jj�:nyeXj�M���+�v�5�y~����{�����,8`��j����b(�g�|_�"�7\N�|/k���Sw�⑓^�[���W��snTN�:�Q��S��Y�,'?��H�M��=9>����l��&�L�FJ�3��)��ʊ4&+���f3֎�N˿LA�0<\z��0�>-����L�&��KߚP+�0�˰Ņ��X�_
tj��.����9@���/_�ʧl&��
\�;�X�"�#��j���p��aJ�9 �`�1����j��22���KȮ9���Oq�=�s����V��^��r����z��g��c�� �'��U�����mH^�����l��Z��#�|�-�'7����n)u��U�Cr��q�;��f����k�NNe�8��<]��6�����t0q����:�C�76͵���l�+�h���/Yu��oɃ�V����'���N�4 Qcb�\=%yf�s�-&|���<㭷��M|&5U�<�\�م�nz{!�����	ؾ%�C��A �&|���c���a���˙I4:2�U��RC����	۝��aU��MZ���@d�zY����22���*|��T�t�m�=|L�OӞS�%W����E�J���&g��s��{�񬇒8E3���F7y*��|4�,F�d]��AMނ�y�9(������2N5wM�:Jx7C�|�4�B����+n�K;�ѡ6��0��dԾ�CIR��񈨞o����6o2T\%&=W�h��ͥ.b��B73�1+?D�ƍ�{��B<߇:�!����{6��6��/QiWw�:T]����ֺVI��a��rR��N�}U[���TT!�l���+pcI�&���K�؆7蔅�)�t[f��,]����Լ96Z01�_��t���6���io��9���X^���4Bgæ���(���1�w�`~Ω_�M��Sو�:�#8x`��жW﷋�"I������*����c;�N�+`PgUp�?9�(]����r�$8�(���,g�Ҥ,��FD(��"n�R���Kc��3��A$���d2Ȏ?�n��$�W�u�+7t)�E&�@=�3G=;��O�MX%x�S2�� ܿD�d�l��-��x�� �y���j��I/�.*���(S�
g�g�/4 <�g����z��p�i�B��@]�J�:2q.-��tޏ�L��ɮ��A�ο�u��LM]�h�<�7w$;`�e��\{��ܧ�G����y�Q2C��*3�D���œ��bԧ:��:2V� �sy���vfu����kڂ�4�c\qӞV�Sش~�[�� �8 ld���X����H�'#!���J�7��?N��ό�A����3_-pI7r�҇O��h�om�\
%B �A�+�?%.���]���N�N���2�>�����dپ�"���v��q��Y{�8��ZbF����WI$k(�c�yt���N�S�{�{��23�~������y��6}}�|P-�c���d�D�G٩���و"��BD�5K K��V�*Y4d{���4ȿuE��%&�8i�A��q�e��IH��?�+���V�E�[*3/��{��n����kɝ��˦'K�oΚs�r�l+���8����5OUrIdg�T﫼��@;��G���\_�L��W+E�:�}� h�"K�?7Dձn���/�CU��1R�f��8<�+��|.����m��D�k�-o|�@�w��3��Y��E��'�`�P��(���P�.��)z `9��e�+�!�*$EtO�����}�����SF1��Q]��±����s��ߡޒIo`
&�Ƣ�'�l��o��8B�e��g���/8���7��[�=/l�>�-�ş�!ܝBG��׼�{�"����c�ޏ!o�˒Q��e�����D�	�+KXpK���o���Q�oX K�-��j��I�O>����B�4k�k�+_���.ވ�����O�?�hf��{ȑ;��\̓8ƪv
|��{6�I�*�O�mw楌�ykeĝFO��:��� TL��m�)"��������S�U��� 8D�Xv��]Gp��N��=<�����!E������	#S��N�}�ه�q<�$N������b �#Bh�&_{�������m��Q�h����hiKN͆��ѫ"g�;��U�x��ɴ��a�d���Ӡj�4k/�(e��^�r�zM�z z��.�uJ�$C���ڙ��-�e[*W��d���F��>���|(��{<�R�E�$?u!EA�K�W�qg{�����$q��,�#����(c����B/������	
�R3AkBL3?0�,���*O�ƫL���g�JUA(v�l(� F3hT����}�/~�k��9^*��h�#Q{��>H������>#�cdh����7���7.�;��!�m�?RΦ����-���F)�V�"�	!,�w�)Q>�!ia�� �����{���-b}��K�!��vw���*I��Xt����R���u��;��ܘ}]�Z���[��q�k�c���6hOzWS�|e�P&���Ǧ$��_�G���G|�^Kf�UT��v���Igi�m��)*�zc�[��J�G����!m�L��śoW��XRr���"�s������ţY돃=��9l�[ƥ9eTٝ3�:Jr"�h�N��4 }�m�Jf[�2$Ѱ�%�UM����-��Y�׀guB.�l�/~O�R'N�������I�:t~x	V.n�z
���LV�?(&�vξ��0˖8��x�(���o�E�$��l��o:g�:�;�R��F�"9�L>X��Y� �I����O��
�h"[�����b�b�8�L��K[2�'������+Wd�B|�q1�!*����p�+��^�?c��6@���&Os�Ý��2����S���@t�:wimw�c5��I��-��Jv�>���s�����r�ƫ-פ$��]�������Lݣ�ce����ҨF�½�}�A²y�!�ٰ�=���މg7*�J�N��"�	~ۣ���B��_"����_��b�7~
׃�A�V�)&~�ÉoC�Af��*~ue�
�sm��&���D�>�r�
ҧ�=ov6�&{Ɏ��!e�;���(ׯ����U�դ��p+�{Uj���-��J��4WH珺ER�	���Օ��TH $�3�HHL�mֵ��Y���=��A>ڰN<�wk.�D��IjT�Y�~��X��"���+�X��g����
��\3[V^�==���9)�o&�&g-]r�i6�|�y�n��lF_����8(�u�H
 2*+�iDQ��o0תI��n�2�^� ɋ��J���E�G,��I\N�$-#�wDf�S`E��'�id�ޮx�/�����ur�JH��w}U��J}}`�ü��SD�ְ�rR��7wرb)ְ�36�"p��Fh`�[�2�-��L��w0�%���'+���-$s����]C�s�'�PQ�/L���F-��*H�衚���H7k���Q��a�$�"�Dܴ�����s�K6 O�,̞�}#u�m�j��m���4��LOY�U�:
<�/�5}X�,'FuL�Y��t(����8�JX/���@U�Kb�'�J����d����sT����H���$.�wn�K���y2
�m}�QTE� e :�~7kD����5��}D��Bۄ��Z	ey�ЁH�P���SR����w���o-`.�Xt����+>~���6y�S�n����j5>�
�������*ð%��S�E%6����A�`���ztL��g�����%���wVH��}��+š�<�,��Y����+6�KM|&.cOyP���ԓJU�7�d,���!z�L>jM�o^5h�;ۖ w� �����,���
�i�v0ɛ�Tx:9��Qb|q>T/����[hѾt��bݸ�.�C����Mu@A
�^�U���Z<�Ft�o�U2���⛎��k�yV���O���qu�a��b�En�}�:a��94� ����-
�̨�_�η]I/���`������f�δ��p�h~m�rZ�@	�f��+�~�B��~Kf �jmlةq�l�L�nf�����2;ǼѻN
Z(�	�O��A`I.
;��������+�	�J$� �tS��GO���:��xF�L��2����ԏA�(��L~ݭV���Aw�}��[E,�q*0�Е�� ;�����)�K�v^/�57W�ժ
p��]�6$x�n�#�����a�V��v�7ř��QG�d��b%���q V$�4(���(l��!�P?����]��rb6��;{M&��IwMXR�JOhon9��>uA��U�޿Q~w�r���e�x~����w��/��\+���f-eQ�$�����}|��(8�\<\ݘ̈́|~V���٣����PeA��c�[�p�3�<��CxBW�r�㗆6��%B��=�����ͤ/N���4f���ƔLW*y�!��K���=9�A߱��M��z䦑�g�"����&��i6���Fo@��l4���9ٵ�5Qf�g1��f)eJ(��FJ��r>ɣ\��`1��,X1�(��p���Pz�I�?�]�+�g��G��l`���&�{37�Mg/"�Ed�vP��B���k؏P��R��f����M ��^�?L��_p��N9�y�t~�z�EB7��C�$�ⷖK���=�i]b�|ʷ�|s�Xd\NcKQ,�tU�"�Xd��.�qK.�������WR�]�#��/����Ӧ��ez��ݔXi^z55�W�C{��¸����!�|�|��,ع1~�$�x"kë1Y!K��u���p�
�@֬q�-��	��O��)�������j^�_$���s��� ��D٘���ֆ�&p�J��a���t}��}j�t��Pnt!@��_��ȥR�k1_��=�M�qY����<�뉡�M���yA�������Cdz%��mi%�e;����W����\�c�P]Ԋ��"
���z���z��	��y�Ѭ��b�6�[�j�q-�^�	<(U9=g���RIRG�H�<������u��ݜ��c�7���`aY٬��ҮlU,C�&����!���Z��ޏT�� �`�?�!kO�/�q�3_Ū�}_�:X�q)+n��!�2��^��y�����	Fc�u�x�#2/)�FӨLu������zH��(�T;!��"+�%�I�k�4�Y����r�,�B	L�c۵(��G7<�H㓩�\�J��>Ґ%)��ux
�f�+���m/,����v�_�!�ф�?�lg֋��^�Z� 5W�xh��/�("Υ�P�Rv��CP�(�Aj;D��R#������g�o�j��ػ�8�k�<y=��GwWb���i�U� -p#�:���UGֺYӨ���R1��2}�g+D;j?s�؎(��H%wi�`���x�v��� 3�Z�}���?i�^�2F�F�	�/���n<�y���3�Śc,�&%�"ok�#@��:�W>�'���x{,���Bu��}K���/"S���J!���S��n�rC��ꂷɢ���Lȋ��GΒ 3�."_�F�D�Z��=��kiS|c��?�u��G6J�����2��N-c��zC�2`�ūa]#�������\��g��=�*�"#q±~��YFֵgQP/���h�����4�^�¾MJy�Jً��Vڕ��x
脮��YŴ���Xp�����ft�~l��F�l6���3�3;�+5���Y��t��*Q,@�V�@��U�fD��}f�N��h ۛ��_[�>V��=K���">��R����'}��N�"3.ɳ�0u۫~�rv����O]Ggݪw�x&�����%�u�Cl;�#ȤX-Tj�Ռ���)�e��!R��r%G�T����N���e��A"`���&�')�e1�����)I�B7����b�C�JyY���e?*�G"�U�@��?�D��1��c'Q�Yj��]�cd6�L������mۇ�Cz���y*w�v��`��6*
Y�������(/)��љB��R�f����݆M�D8�a><iN>(�b�Ȧ'\��$B5��}�$��YHQsdI=e:����u�|�?��shGx�;@?ĺ�)1b�g��}�.3����n���ˣs/�2CZωj��I����C��"��~[�i�3��	��e�R�� ��g����_?�#�󈣛�`ƥ7�)��Ҝ*�*ˡ�������uㅲz
�'ϣÆ�PK���`�����-Nj�،�B/���#0¯x���Id�3kW��}P��)��b�"=;�9�/+6qxs�Rg��pK/���;Ȯ�8�m�zBe[��c?�� �3�X����jUy��q2O"">p��9߂�[-�v�s�?��r7	MiG���3���S�y�\@s-�$8�+�µ;+�R�
50y���)��ۙ�J�����_�R���U\u�.� ��a�F %�,Ρ���Eǉ�/���Iߨ�Ւ��K���CS�����o�ĨI�I|�{�'_&�2��J�k+[���yҦ����Em�bz��L�uh��rz�6+�av^3
6奆�磯�r��5z
���-<�0eB����\��g
�+�AW��O=��=�e>��>��=�p���ש>Ƽ�t(ї��usWg\bw@�~��(��Z�m�M�z�d���14�?Dsݴ�?W�����啃d>T��5�b�I�;�,��}t� �1�Ł��_�l�����u�<��
�p��e>
�-����=B�dx�u,�uA3h��ֱ5	��+1PŎ�S��j+ۦ7���Z�S���&��f��%	B�a;�we���p����׸��8�[|�F�O�K /�mm|P��Ԓe����`�Ǝ>�p�����T͉�>�ɔ�2|��J��H�YD�&�H`�T��2]{�����"Q3�@�~;�`3�-ͫ� /bE`��B�!��V�8ľr����E����<x�<��%g�b����C�j��멊���iʻkcE�t����N]M��JJ������"5���"�[�B�ܲj�4[�&\�{}y�aA(Gk���]%{�=�%3��AۗHzyߚ��w���ꔺ��-�Z&���C� �g�����V��������|!����lmj������%��
��Z�(b��k��G;�=g@B�0L��oX���HK�Gv�4�P���Ld��0iOt/)y�`�Ɨ�'!P�whz�v�ss�㘆A���6!�1�1�M�����K�����q�b���U4�Gͬ����$П�I�m�{��x�-���=g/�������F8?Ү�z��W](��S�K����e���m� �ʎH���~u�Е�)ȷI�E�L��*�D|o ȕ
ӂ�c��4������f��~�"*�\�M]v�k��"-ҳ�^������s��X��y�Y�k	 ��?��ؖ��֝�����.����,N���+O������s�ح=?G��K�x1��m~zA�5��IT�ǻ����X. ��+`T�< \4�-CT�"̠	�8� �Y����]��WMM�S��`�	(@1|V���
����!(����*@�T���0wk��P<��*e�b�RmjX���\��۾Ӷj�0Q������"���R�i Xoi���@���i|��YQ�79b�6bu��r��tK6ԟ���nuy �E8�C�F��)�J��Pax ӥ"�+�����Z���:��~?��UѬ�^��9=I{ #���jҒ�"������@��Z5�9�K����=��r��K5�nH���Rb�K_~��XF������ȶ[��m��������u���u���� �=��IvHG�²]�k��.I�� �U��y7
�쨾��Y!��
�3�<o�Ĥ򜐊�V�8f��J���W�?��B�Sg���gEy��B�ǣ�
aD��xN���������K���B�X�t�=g�k� 9��$�,���_��l����I�Ԉ��G
����\�xl�����&�>�mUYsW�!��W�$P5�^"C֞Jۂ�+�qL�l"hs}cGnl�d$��z���q�v3��7��ҙ�qi�2�]��5�p���@��ړ�F��j�	��V�4K(HSe�Lx4=Q! !#���&$���ϡ�����
����*q�W���Bj����"�H�G�+�j���+�_�s��4FE	�w�oz�B�ZnP@<�^C�{�N�嚊�ˑ�Gp��I��_L���c���i�	`iA��Q��|��A�+\�ۛIvr������~7��99Fmo8H})�A���C��99��M�Miֻ=���z%��8�����s�&?0ݬ9ӧ��W�׿+^��w�B�A�(4p~E��H��ӷ�>���U�o%�i�-vc�Lt�+��ǯ����s�1s�;ǖX�|�_7J*���E>d���ُ�	wb��NJ����?*�8��!�c൓v�� 	P�0�pQ%��C ���*�����GK}�+�=��ls��Y�&N5��㭆��M�V&��)B�V����ޏ�� �	�+ؓ*����w��(��M��i�A@���q3��&�����GMo��X���7Cn@��

I9hP��+)[ 0[��1�$jA���[��`ӹ^Jw�*���Pi/Y�����W������D����n5�JN�P?��H����G�H�N� �cf�(��~���]��Z/(BXci�����%y�&��@_C���~*Kkf�Zh���3jZp�A�[/+n�*7Z�W��#:TYc^ْM	�#F׳�
;[	 9�O���פ��a�
���|�dj��su���i�>�'5�9��~4n���'��P[ڦ6�2_q7ˑ���R�}p�bG4]�j�;�Î�� -�t/v:\jh� O�-6f,���~d�xO�r����ao�rb]����t���|-�۱�ɨ!(��b���(��U
��4�o�����Lc��E��e���	}�=�řB���[ڼ��j�	B�8k� :��:P�]��~�ِ ���h��{�e[���y��Vr���b咗�CP��
/3X�����
�/�C�t���9k1:NY	pI�P�M=!5���S�W ���m;��h�����R����v� ���쏕o�ՠ3#_=N��l=	E�}�+{�2��&s�Ks�m��"rr;ݜ�@J#۟�� +���o���@-��'�����L9�'��ͭ��V��m~6���ψ#��Q;y�rh(ފ��w�2�Q?�F�;5���j�V73ㅬ7���q�oh\�&Z��BY��P��f�d�	y���8���KфبK���Kp; v�2���L����(��*�D@�q�B|U"��챽�s@��<O@1�a!'����ѿ-��ō���K��(x��wyK�4
9,T�&�	��7�ٶ]��
b����qmacpP�\��[	0Nk�3a�4Z�?rz{b:o%�:�*��-
B� ��)2ZBp�֯�V�A����2�Xf��HO�l)d!�N4V`�Q�lv����7?�8���L��/�~4��Q�R�wiǭvQ@��9w�JT����-��E��>��(^|�Ͱ��~jу
M��@��XwǑ�s�*��M�l��on�V�1b�LT��1�*��I�/��&�=��.�O�G����	��Y�b.р+�x�Y���M�g�Ace�W,��-,�#�b&��xkP_k�%s릛	WOIf�蠢�=$v�3���:���@�ʳw��=2����1bn>�"kaC��l�_I��X���cP�	B8N�Ǫ)�ܶ�7 jY��3u�ywN��"8�����L��'*<[濟H~�E����Ѝ�ݛ^ý�"��K���>"l��RT��g8�QY����6�J����%�Ms��l9�O	�H/�y�Ԡ:�)5d�@�U�m�:6���z�)���'����/�=���"q��˳�焆�; vұlsR�*�O ̶�k����*�Y?��4�XY<�����[�\��M�*�aW�ↆ :��v�7Pf�&�;s��\5���� _���7�6�Ƭ�k���	�+:�w��Rl��#x�TJ��9���u�-|K�[n�f�I��Mz@W�D���a���[]!��CbD�j� �u|������X�7�S���2�PF���<���ƈ�ޚ]F̃@�*����.���ɢ���U���h�	�%|Q�(��n�uN����
ZD�V��+�=7l�f��B��an���t����bz�9�>�}A��1Dbpx�������%�u�4^��U�ԋc<9���k5��hl����'m�Y�݋��\��n8�����`/)�"ū�7:��S;��T��R�}n+����2�4R=�=z%8a�
�nǁ�֛���:a��08���z��@eX}H8Pb��aO��8ʂ����ء��,#�6ہ8�$���-Rh
�G��AK]mc��/�$�eZd�_�΅�ud`6 0��!N�r!��=�ݙt�1�|���9%���?���P��oZā8i@�g� w^����r����O�`S`�����zA��"�5�Yg���K�d�R�"yŤ�*[�������<3�]�Ŝo�Հū�c��R�nY*��d0[�q	^&I��_�Cυ�q�ė���ۆ��8�u5pga~��N���4�	�8d*y�� _�Ă�(-N�ݴa�5q�:��aO�a�l�9��&!�iŋ:ȴ��E1MH-�K�����V��ш��ȢKZn�0*�kh5��?���F!�����E������b6�����T�n͒Rk@�-���C}��[sr���=�!�S���"�0�2��
��E���~���C'-M�4�|#yV.�U��zټ�� �m�!/�!����\W�O)�9N^���2��6��EY����P��q�7i�PǲҜN�*��{P�W���w��@�f��Rg�M�\�F�突*�U�Z1su	_�l\y@H�W|�w86��������%���4���0 nI����J҇��av�Uu�*�_ۃ�a(#5;}䝚%����qH��ת��{�p�����0���%Rׁ%/.D�Hr�^"��@Y�7^���o���6pR�۔#~Ye;	���y�����ը�t�D�-�!p��f>F�5���H�jP H�iȁ���)���!	"
W�k��}�
i�%�%1VD�n���5e�TC`�ީ8�}7�o�{+S��RLa>1�A<̕��vE�2R��&~u'�x�j��S*���E�_�������WS��Q��&)E��dHF�����l@�	Az��)7�$�s�����<�')�4nx��'Z�S��ZJ����j1/���ۻQ�CS�|/��oR�T���+��'�
��W�M��)C,峬<T�f��>@��ň�虼�'QG��dY���3~I��=d\�/%�j��w��v/��<���I$I-A͌S�	��<4����'{�8��9�ٶ�ˍx��z�b�pWbի!v%ؤ9��.����ZD�L�"u��"��7��3�\�R��1��
4�[a�,��_�&���p��}r��N��!4p�%hC�f�J�0<�Gx�`W�9Ng��.JC��x��*��/�c�Dɼ�ګ�,�hiQ�uN���;�)��&=[>{\��X�a<��,HY2�o�W���nm5~Ց|$�N�iЙ#��Ij'B���0�B�Z��}�,���%����N��-n�r]yϫ���54�D�T�b������!����U�go+'s� � ������/�������Ї�*�d�r2����ů_	�x�N�ģf���1J����`RF,(T)� ��E��ѳ����zK��<�{����3��	�&1t�M��K���������P�s:�n��kL��eH�q�.�6s��J�ĖJ�8�T���?�Ս� G���R2n�_)�k<"y��) ����eW!봟�e�k�kP�=�?��/	5������WJ��'�l�A)<���y+iu��tv=�`� �?$L~@�u��y(�0��	.����	�$O�Z�0��|"�����FB�!)��{e�^e�.g5�*�7��m��}d(�Zl8�i�s?����g�Ǚ�}�j���m�hp+R��JM��q0��E��䜪��H)0��R�kg��l�m�u� ����L�<e�,��Y��������l:�mD�z��9.�_I�SMz�<aK�v!k<��%�R�F�o(x`�K�޿\��@���R
uT<�x�Z�hhE��w�x�z�%�����]g�G>�=2�z�ҳ��w,-�/��;�y����L�o�S^�!�$z5��v�L��:M=B��l�����Wy�����0��I�!A6��9 ���fx�����㢧��wv������ݸ��A�Dx���%s���W�0*����Q���zz|&��U���5J�+8���0jp�����T]� wiJ�,�z���3��3�dwQ��~J�r��{:#u'� p��~
��?�PzU0Vpn�v��KTv��<�BT���T-7;�k��/Af���9�$���� 34�?��������d�D�-(3}�2v7��hq��
_�hS�N3tߦ��rͲ��R�J�%t�x.���H�����������K�T|�1�4�]qtʶ�tm��]�D��R�O�{�p��AL���O}MA�l��ã��:�v�C�lيy_(�aW�5�􃒒�L�N���M����#�x/k�>�TO&����疇�5����[.���\�H�%�T�w1�֍-F�%A�m�`��i��]f�
���$���t�w�SKl��!w�U�6�&C"�KMYƙ��A�k��ʹ������TV��ۑa/�����>B7٣Ҕ.�Vy)'�!o ��Ľtǲ�~\j��&��p�$��#4z�p�x]L�\޸�K6<v�L�2��A6|*5Tr���YE�+�0򗒨� �^=�t�.Ƭd��I��w���|��9�t�N�*v�k�ũI��d��3�����g�����<h�g�f|���[���#������3_(ſ��n�3�߮=���L�42WR:c�~�ߪ"�+X|T�	�F�)Ќ��3~Ɵ��+�D�����ɵe�4�\g"H���7��FW���'�Q�P�����<��5�CsQ�w�f
kc%�*T(m~HwA�	V	8&6�����"[qN��p�sBbNH���k� �検���"��h��(����Q�V�O.yn2�rsŴƻ�{z��wn���G2����(�`B���+�O�]���~�
G.8�	�:���J@7`���T�p(�x��R���Fڽ\cy�.�yV��X�*��06H�����;�)r��a\S#/��P�C/��۞Һ4&2=T@���(�lq�w���Hٚ�).��W����� ��U��?x��Z��(��)	ם֯`s�	9-x����}���{m�o:�ga�����%�������D����Z�X>����亗��5��[	�yE���{A�70�&V�z�ڜ�x�x����V�D.�?8p��cѮ2�5��MM�����P�e��&Dy�䉥׏�·�P{#lA	������{���$;�����S�vRY��!�cw�<��aĊ69t����	8z������䥼�swr�e1����<�%>n��ur�J�A��d�6�?���+鍶4!��ݗ1�,��	�@߾P��W��т��61	�9v�0�< �=�n�_)��dM��R�][�t��Ç]j�.�ݞ�k�s+�/+8HP)H`-Dv�q�(\��e+p���%���������;M�W����&%=G^q�H6&&Z���@����(��T��R���0އ���t*�xb�T\辮p�"�ۧឥ�
�1IaJ��ә5�Y���}������T�b���:�Ԣ{%3�2��TŪ�ޥd�2X���kle7�S큨�}�1O��jq9�\�讬\[Ji"��̐!ȑ��z��y&���r�n�?e��5y�E���q@���A8�C�B{�3�H�֙�g���+��\L6��Ge��:R�A���p2��W��U��wp�"����'يMt�!������r��1	��thS���'˵q��J�ʵ�9��t�WN{_�t����E�3�n���G�O�ޟН6@n}����E�h�1�G�A�w��""0x�\�T¦��	k~C?��N��sԨk+1c�3 ѲE7F��
�鶾�Hᦞ����F'�l~�ne;�i�I� ���$�X��Q27弐�4t6ns�e����WFE},3�d�[a$�ހ0��8 O��*W50���N�Zo�3@�r.Խ4x,<�d�J�\����Kdc��Ӭ�Mji��T�3�!��@:������+��/4+4��2m"��QF�B�x�b�(���>��Q[Pof�2�Ѳ�a+������g�K�P���@�ʗ���y�Y��'�PG�t�d����e��_FЊ� ��N�GsM��}�O��K}Ѧb�#b��{9�$"m�/PsOb��/�C�����O���}�sj�Bh/���ku�=ƍ�a�'�DY&����"���r����1�@�#�zϯ[��I2p1���?�#P�����	���w��1lU� 2l�>�J�zE�i�܊ǒ2�N�{��uo��Z8l��|�=��;�ܛiֵ�G?@mo�G�[��g�P�ۑC����cC���A�O�_�1���<IZ���94�Y��i����$���}��5�c��6�%7�B-�]���]H8�$Ԏy2�T��v��EL������F��e���\-,���r�8����^wu��6\Htx�!�W�4s3�6#]䑁����4�
�Ԓ���{:�q��l�$�V�(��b�q����>|5{��;�$�6b�K��b�D�R2!�M=�p6L�^��8F���eG��g�7�i�����J�����AY��B�sR���`U1`��w�N�R�aHx]|���J�N�����s��Q���u)l]�~��SE��Tǘ]<����49��qlG
��6�v�o�Z�
8�9��䠚^3Z=@ݿ��t遙U'�GW(��}�}�~�Yk��̌��Y=b)�C˰'��%�gU� �٪����fE�w�T��3e���1dm����c[}OX���k��d�	�S�.����X�L;�
�f�k���##s�aAq��[�zY��.�������򅽀-��Mu�5LR<�����?� \�Ȇ�	�����]L�܍OuT�s�F�hE���x��wc\L�?q���B��m��L�08"����햠�L��L�ݺ�$��Ӫ������+��r�uC��'��釷!
9(���U�g�}'��rzY����.D��h�(�E��̬&�pU�'���`����}����żxQ��Q5M�����1�O��3Ω�G����P�p�� W6޶���Ӫ_���ǲ+���m�Kh��*>���Y�#�q�n�rCY�8�.�o�|�A�^�"t�mz�FC�~F�P�Wq?O9�L?h "�GɀS���%x��ը�
�����;�������R煛!���?k�i4%F�_p���gsz��T��E�j�`�*0&���+x23WWs[*T�hl�'�E��{t�4�-��{y""�����	~�vY`��-�%D#6��X}��)����w]�okS˕�M ��	y@
g�����<Ʊ��t:�.9�V�'ͻ���'�9��n��ta���X�0��)�8܇�I�J.��iQ;���+���0���z&@)���zM��)?plP*"�_]����ן��ݬ1�i�����ZF\4/?.`2�4�ԛG��d��Dm&�dTƆ���!��ʝX��&�z�0�����v���)����)�)o�ۖh�
�T)��y���>�"�{�}�?�	�G*V�bl�0�rw'�њ�lQ\VS�1U���헕e&���CR�f�kЅg��������oK�/�=ѣ�p�rKW���'Q�e��d� +g�Ք��Z��2W����YR�v$�0�V'e�����
�X{�|�^�԰Zryne'�~:��קpr�?KӶ���r����G?C=�.��*��Oh���h(�7�� ��?���抩 �6ʫ�s̝�̤�Q6��Y��mݯ�Z`��K�F߽ʂ����8��@͢�d�V��76<)������Q ��L���ȭ/��W���R�!7ˌ���D���-�_�X�&��	�Ҽ�2��+H��2����I��(+�Ӏ���g��$+�k�sC@�}��.&�p6�+<�C-l�(+u{����tbwa������)r�>~�6������&*�}JB4�kTxוkК���n���+\��p�=�c��Z���� �.j<�a ��df�ZlI&�F��q�����C�܌��©{dʃ/�y�AP��6X�����3ke(`L�%ٹ�V�R�*�a�v�[��݃����A~�Ҷ��!:�A��qZB������6���[�.[�1�h.��k���["���4��Q!�������Q� H���]�1��.�d&����I#:���/A��d�j��_u�s<W��3�M�ٔs;�o���}�m�
9j�qǾxvͰ�Ӂ�8�v
ҍ���
�jܺ+�C�,q(u<��i�����D����o}򲩹}��G�F�����T����}��!q�3�x������8Ԝ7�gЛt]��Y<݁�z��2(����T؝��j�K��O�K]��k�� 
Qӫ��R79��
*`����T��젙��(re��Y�������Qr�µ�1�ص0v=�t)���G.��Q����'��S��W6F�l���5����x+�k�u��#e�҈+M&~Q$
@�y��?�e�3b�;s��DP��;�Rw����8�Xv���|��ۇ�`+���i����N�U�WdM�Q;2�1���4'Ut�!��\7k*� �C-]F�|���%�YKig�#���u� y5���@fk�Үs�Y!����ó��LE�jFR8�͈$��w0���cҀ�*�JR,$���V����}����.3�Ȅ�eNi�	�:�[ˍ�o/��9��R�S}�F⨝Ka��y���k�晈��@؁i�C��q���q2��mؓ�S�a��S�+���R��Uf'Sa�S67��MW��GNwŤ��)Nf�X��}F����\���u	U���j��Z&�F9^2��<�2m�h{�?"���8'QG_� ���D�Q� [����>qE_P!/ �	�aՇ�V�;*w���,�U��zC@Ko�)�%����ј�r9��f��~��2yNЊbڛ�D�N�<�X�tM�������iX�r��ґŘߢ�E�8%�N�Mn3�L��EO��$醓5�%��o�)=c��0���Q�Ԏ=�k�̮�y� ^�Ā30�˹�Vu�SLW~#���qk|^������Aw��ce�J�p��N�X�/S��J�KrH���>��/�]#b����8C����l�)y�ṱ��l���\;�����
����(9��M;�gQ�AH���"'�y�L�Fb�:o���
��u5Q���ljP��Nj(2�ТtP��'vxj��eܧ}+38iu*�.+i/V\m{Qz0�/������c������T���x��X��P�7�=Ho�J���[wƗy�p�Nm� ���[��8xD_��ڗ�>ct�4hR��*�8��|�[�Ϙ�?��;\?`���L0��S�[#EG��K�~�ɒԹ=ٷ{4s�@6��،�M;����u	b7��WAhm_Y�p��v�!���6¡o��0�P�S#roc�|�i�˦EK����LT��ic��^6�7�쫿���=ؤ4�9͑C��R��A���I��:a폚DP����̈��/�<|�@�����w<��G$R͢�LEړ��3V���� jP2�x����b2��=�i��Zl<1�M�F��S�]�
��! �:�v�0�w���vL�]�^74�/�E�9�В��.N8>	�l �#��>O�ԉ�o>(�So�'o���'�j+���N�e�R��~'n�޶%���/�����n=������`z�Qq���@�^~�f�GF��j�s�@H��=+��І�P��Z��Co;|lJQ1-�5b�6�Z��m��.k=����E*E(��/!;K����-�}������v ���b	�d��ˊ����$FK�؊R̀�
ztԞH;
�m+o��ilo��T�n��|�J�G�Lzpqf���bǏM��b���D�x��-��o�5�e����~q�7v��O��<�i��!/���ui�X�3���ɩ+cgU�pMB�>-��A+�s�2X���� c㲱*�kP���:�j�	Y�N�5�`f��%��ѴV����y>6���Z"%A~r0��k� u�����s�t ��πRښ��N������Wa�8����P@�wd��I���	'�Ӑ�Y��6U��_��˘|��'��1V�4�I�ff;�"� j�p��F֐eNtDyQ]�t��iO�'͈�=6�Z���,qq�>�l��,����f`_�dP�v��w�T�4�I�D!���b�~�7�?����B�l��.lsب҅b��-���НKGh�C^R|	6��`�aB[���C�>�2o�h��"9��cB97t�V���sb�ut�}�l_P���vg�g���nF����Lp��
�l#���yRJr���}�1̴j�7�:T��9<�Rq^C�[�ߎ��'#��n�C���/���BT�Z�ҥ,�sj�m��`��4nT7@:9b8vJ�v�܎��% ʧ_'֍�Hn���g>���+N�@�Շ(w�ƍ[����.HVN��O�倜�r�_��w���l�c �yD�h�ȫ���`&<P;��vd@�^���Z_� �Jro{p~�piO�=�q���ԕX����Q��Nރ��"���%�գIܒgJvLA��v�Ft,1%����B�BS񒌗���h���1!�|�/��v��L��A|ghdw��_�#GQ@� ���[����_�=�{ǰpMnY��*��0��Z��>��&�	�}v��Mh<��ye�`�l�i�S�Po�y�d�̐�OCM7��SR_�����H��ɥ]�R���{D���gA���;�A#�����-Y�������V ��ʉ)jSS�Uvq��7U�]��7�D#��"B��T� ��K4�i��"ʜ���1T԰�1��G$��yEg�
����
��DT4� 0UA�o֚J�z����&�l���rp9��Pw��BᦰT<;$�T�r�"x��Wj�)��J�m��O�u"�,0�	D,1V�d$�w�Ű� �l�:�h�F_2O!3�}�mV��h/����C��.tqtgu�訚�&�$��cO҉��,?��`J�� �|���Yk�����@�J��
��g��չ�AyxY����"({���4��$�jڞ~^En Y}޴D��u�:�%AXQٹkJ[��^2�}�3$�b�����˕����Fk��@��hq���ˍ��pj�yp*Fn������S2�H�q��tji�-��t�D2�VV�B�5:��"��� U�e�L{����������:%�vn���Z6s�՛���8C�%,\%���Y{�G�@�ě� +_���e��7��{�'kQ&ͼD����@������F����a Q��H�~`���f^U���� *k/	U映+M�
wM:���ȷoϩpf��o�Zc^�h��3��<dxGῖ�)�L3�^��ȧ�|C�ɋ���jg�U�<��?M*�L���"�0�V#,��>&��;l!h��n�Ы��� 0nI��ԝ�E�3�(F<��OU[����ݗW+C���=w�V�J���#�hn�h�M�\�[�H�zni+9��Y�r�뫘ᕉS:�-/�� ��b���&����+nmh@"�in��կl��Ɏ�7Q$Kd��_�=�(��9��)��=%g����O�B�o*��;^4��׉�ǜ""<ms UYJ���=N�"�v�b����?�Δ|_�����=�G��kՕ:�Bm_w6�8�	�	��%�P�
��2b���qO32̰Rzn��Fm#ܵ���ɝQ��L�W2U�q��pϯ.���.�,�Ƭ�A�e��Hnwk_n+ŗ⊄�ݣ��֟B���Y5.��[�k]4�QL1�:���
��Ų�L�mX��$���AfQ����;�X��Űv-�]y8�P
N�\[���,.t��ֵB�*���2[���h�.ݶ( �fUY��Z71D�K�ӳ���8��*~0�{-��+�^�eH��^���>�n�"m��O� �:󞍮Mj�̂�w�{��Z"����cv�sX}�,+�'Ĥ�ڣ�������D�w^CH��/s��W=�����_�#�fF�!��š�ͽ��M�_L�'�w��	(Ʀ�/n�ڛ�Ce�� ��h��c��({oW�ج��0T��$3n_�L,y\��;�x��Y�5Q������MO�KXb�vr���)�Y�Y$��g�S��`�u���|������.^361�x�W$a3x�ˆ� �V{@�f>�-ڮ[{#q���N1 �g5�Xޕ`D�sݍ�3:��_X���cÒ�HХո�h_-�����z�]G�{+x� ��ˠ���N�j��Rb�i׳��s����z��e� ��77���X����E��Fl�*�[	Z)H�^O>��¬a�"a�t���Y�0�	*e�`�~����f|��"H��}�&H�3�s2�����������n.�/.���d�&��r���4��H��H9<LK� ����-��z�!�&&ິ�G��;-Jϡ%4*�1�E]��} @���n'3rw2c�5��ȩm9����Oŉ�[p�'Qv��Z�{O�l(JH�
Ч'��	��� ��s#��p'*���G��y�&$����Q˵�<ǵ������8N�����iF�5�8�tP&̝��x��	[��
;���PMHII��}��Nh�d��c[<�^q��v�J�\�M/���vI�m)f�%^Jj�MB����������{���L����n�aH5F��v��_�N�|"GP] ��UVw��T5%��E(�L��\ҫT�-�䠲�Qk��R��cމ�� ��{���S5� �l����
 ?���v�Y��gk��yK�������qD�y\N�5�.�ia������)���À(S�8��=\����#��c�����D��3��-	7��r]���Y9��*-ж����$����[�3�R\���53�������B̗�,��P|�IǤ�&��9޸��U������uF�Ķ�qH���t�S�"�����ZY��|D�\̕ȫ��b��+��r��a���2��-�%��d��X���T������ k�?�^^�·�^��C�f��ŗcϟ]qy�e��=K[Mr�x!J=���П{�.!S׃?f_���觨�ё�J(u��#mO�C��l����X*�BN&{QO3�Ŗ�+� �ԩI3d�$�����������
���	���u?~F[X23i/��]������@���MV<�&�=���{v�7�1ڕ>pƊB�\��3+ǯ�Ҧ,����j	����[��%JsT��N��tA0	�8�$j����3{ު��Y�3G	T�\�J��/E
�]�/�@qU3����TxTPY�)$�����T��{�R-�9cA�؄|Յ�<�(m��t��\U#�& �j��k���Mv��� o_C�`�)����mo���:�nqb��a8�:%_�$�Uv~�U&��~#W��{T��v+ݪ��<��&+Jx2�z�oF��ϥ   <q�u�4�Di��=G�0|��n8�ٛ��"|�Vt�@8��jg�Ylڃܩ����� ��ߟ�=>s�NMy�0��W�I���4�P��%!%������1&Tܻ���Y�ּ'���v������^܁r3So�f6��3i g�c�A��N�5W�����NuS����7�Y�]��-���R���;�gI���T�)�2�)/����M�M.���^��,ŏ���� ���X�*�L>#J���f�a{�"Bl�-M��~|#6%���X�?�6����uH�* ��7FU��D�;js���>�$0�'�q�
-�x7zK�Z�9j2C�;5��N.�=I�$�;R��嫕�t�D0�������<�@b��0��C}�wH���Ĝ4���f��)Pw��RF[�{z������f��q�ny�B������ۨt��8�U�\�,��#i����s�9[�����"\A�p���⸷}[㘋B��2��܊��'u-5R�,SqA5P���uk�S������L]Gpƃ^��Zǈ���s46�^�R�g�L��Ѱ(d-]�:�Gܳ?�cEo���QA
�9.��3�#*E'x4�"���	V��rp$��X�����0�7�bF��Vu�ze���t�lmca?9IXU�-�|�@<m�HN���%�����@��H�Nٌ���I@���tτߎH�dZ;���sf5%�uJȁ�/�X�K�B���T��z��~���Gi�p��@�ݳ�͋fAŴ���e����i�J��̣��XO�t���>�gR���7J�V!���/�l���`�&Q+x��Ÿ=(����Gq%G�3�yJ���� �a����sq�l�-ڜj�����0	ǬV3��H��C,R�3�?a3���>�Q+/���VB�*�M8�~�����s�r�"�䐻kĪQKi��D�q����I�)�a�>�������Ε���{@w/���A�lE���8��k.�L/R��g���R������%�e:/���Ʈ�l���`((�E.7����"�A_�.7Ϗ,uW��%Ͳ)W�p�3;���sw�
�nw(e��ĝ��ȁU�``���S�tp4�E@a��~�:�o�HS�,�!t�ڼh�]��T.�[r$� o�����X��/+�٭v�<��?k���V��Ζ��c~� jٞG!h�S����f�/�ޔ��!�E5Kɕ�'ǝja�ӤvdG���}�g:=�#;�~5��Y��/���������6Hwݍ����'�D�Sqx�/*ZYef�F'�t��Y��	n�X��K�Nv���)�n^v�A���P�u�ż��=�w��w�y��#'[�m�Y],LZ��a�y��h�̠ 6#�Ml_N��y�P���Q������q��<ݰX��-?
��r)P(M3���
��B��e�ulns
�5�xy-uL�M�V	���h��g懸���E�1�z�(U��~#_.��BH#��]��O_Œ���_QFT'S�wP;>�����А�?����H�,<���'�`	����ď�R�-��'����y5οqe!��R�h���E"4*�r������#�[yQ���Õ!f��r��y��:bR��<�Z����o����Oa�)�yF:-����ڈ�5�G��hr�	��6�C�m&�͹�!2�3���#��<mt�6��������-@�h�X�t���jT7ap2�:�Nh����AD��v�E[Ϛ9�h��齖�A�T�����l(6�[9�'׃s���Z���{����]~ˮ��k�yĿ�)�R�!͝���A��d������-���6��>�ً(����z���?��k���!��AΉ��ޱm���P�F�/��V<���۬�Jw�!�c����=�`+��^<P2��~�+Q��0;�9�}]��v��4�.��ذ�"n�^���vG6C;�./����]!{N|�##���?ndI�&�0�2��'�ݓ�N*��j�׵�e�뚘�o)EC���D�"ad�9z��!{��9��t��ZƓDD��Zw�rH,:���d�I>�� :VC_B}?���au��3DsQ���c6�l������������h0F��}G�Y���ܻ�4Y���O=[}��+���N=�~j�i��ږ"ʯ�Y���*�V�������� ֭ s���P%숎��dv65����︶R�Ռ��,sV��=��O�F�
����߃3 ��n�TH�,͓+�k��O�]�����=�17���r�0��ؽ�ݡgdUJX�]�R�>�T��?��P�5U�T ��^��%"�$r��/e�xUoᗂ�E�2)o��P0:b��g�ơH�_��O㖧���:��9�5�۾9�,��U�#?\U%B�Π]U
��J5^P�#>��R
�[V�D�A�{��˭�8���B�І���DC;�m�!l.W���i��Hk�b��wj�*�[t�<CM�j
d,��9�q�a�	?ȣ���%�z		������#��n��#֓�}�`�
P��bvt�&}`&���¤~γ$�|]V�)\prz���H��h��9<��4zZ0��cꏀ�N�o`��R��dq��F��WI�p�V�*"!ِ,��P��x9�{,���Z[�Ǭ��n>!\T?亄���9P�ٺݓOjE#م	�Q���Y��`��lK�M�:�F6���0Xl6��#��+�m�"���<�z^��q�]<oC`;Ϣ����*�\Yo>��󱂣m����݀���4��~U���l��;q��D�|�<�SQ���H�	�'?�'�u<��z�ֹ�C�V��H*����:�M%�M��YB�� ax���-��~H0f�	ɗ>w�n4J���g<8�d�|k�ݤ�@Q�̩DD��� �_�g�������|�X����\O�-L�2��1��\4�"5!A�sR��?��EC�����`v�<�ƦW��N��4;6*/5	��2�0Ahy��F�*m'���@�� m�a~�C��.y�$/��NY9�hh�ĊQ�>wYnK�\���^נ>KG?)ef0�`'X�,+���O�D�j�݈c�����o�����,��Rw��>����E��e��L�L��6Jxz
1F=2�B��!��#�4'�Q�@��Rhg����n��v��j�BwYr`�-���� ����wR��fUl=��{�?������[��y!3a=�9��m6��IR��ۍ��NEH��������mP�[�#��A%��6;�WV`b���؜�0�(${c�|����:�7z� '�0'Ύ�!�v%q���\h���u�!�5J)2�
�-�.�oeG�,�����f	�4�I"��b�Qt������K�!�u���+���C�v�$kB�D���T-��9��"�c��PȨ�j����bc�ˮ�W�����#�ݰ�*�MR�=#��p��G4#������}��$�z�OD�����(�9�s!�Ӌ�Q�^��ev�v�.Ny���L0�OQ�)8������i]�$�c��OXL��C���7�q�Ի�m��ʓ(�0�K%v�H��ՕY������!.�����p��_��ϼ(�	�_(Q�3������橋����xo�c|O��c��s�!]3e���\,�,�5r��SR�qq�m�B��4>%22B(+�@U�)��'�q#!G��𾻁��q�Zk*��UX��{H�4,�����t��P�iN��\�N�j]h|��H����*^��<�/c�x��8q>>����ê7F�7!�I.�O���/�.���p���ld�8�?F��9Y�oL������*n�?��'l�CTB�+�d3��Z��qd���W�22j���˗�O_�^-���BK��/oS�)��Q"){A+�%�o˾q[(<�]E �#;x�kD�d����<��]�X���:4�c�I.3�#X��D�tP�7;LF����?�(�6+2z�Fپ�I ��Z���a��+�T�E�ݺ�P4/RF=JA���FJ41��-EjE^Ϲ+������	/�a��1iNuE#D�<U�[���jϒ�O$kҷ�J�PL�_~�"�/�q	�]������.$����d=P��j�LZ�������bkg6���YMk���1�Ō2TLӫf�PA8+D���c.S�ዓ,pY{|��y|U���K��� � `D�n��ȹ�c
�e�xw���Y�
k ��(&9���}6�����5�XжO��Σ� �!=#�������N��ۙ"S�$�'M�H�UӀ����3j�� ]�d�q�f���E�+f�/lۏ}u�p��u��!�y!u=I��*�0gdȠ�i��|nv���d�%����n�5g��:��9��fr	�y{�\6�ULi\P鉉�vYv�,� q�9�T��n���پ�����.�.��9��uLr�SI�Xct��%�����2N/G�p�dRR.Y�_��M�P����9r���o�@��^������U�kd��=,h�OF�ɵ�$�5t�4x>�8{�JoMT�з&ޤ�3O�X�Ke�^�;R_�}:�?��y}�O��h��*��$ءjb����y�l��6���������"@�;�4ɽC
��-��VBD�(�C��:_���jq⾇z�> ����2�����u�d4�)�1H�E����d��m�����͏�P9Q���<��z��00��+����3q�Ҽꥆ�ݰj�3�1�eqїx�� f2a��[�Y�:r�Z�NUE?mH�:q�<@z�G�����J��fi��x2����j_���KO2o��!Dd��Y�n?���r�7�>�5��$�h�N�Y�!��xj[@�ԥ��_B��{������Z��*l�~#H�xU$L4�pS�9�,���Ke��'�w��(e��BN�ñ�M��Of/��o��k�~��B��\�.p�&�Q��7����&�L :�ۻ\��ӂ�$�2�he��dL�|�%�J��(�2���'7�����S62[?�1`�&/�(��|4�q_YV�ə���z�	�4ۓ�&��L�|��-
�{v���!6� �Ȥ��l����aP�!�0�l��_X���=�0e?���4�T��@o�W�����?��ɵٜ�ʛ'k���$�W۹6Q�F�F�0��SMȜ18�+��{��n.��&�����ZR��ַ�E�|�l{v2$�HK��Ҿ�&d���T %�)5� �?��%�&1A$Q��	�����?�G�%���� �`Y����y��7�ő��Y�O��s{�d���HS4��}n�N���6�T�O"��B����PN:�aRYh���з�́�imiO-�JC/�Q hr�B�q~}���@ 	&G�����!�������|f��O�M����a�baW�1��sthG@�r{��>Ί6ow��T��(�ΘT��X^�6D�PĽ1��.�n�
蚰��� �!���U�ϓ��[*e]�lZ���?{k��/jp�D�释6J�|��q�`� �r�}�#LW}�M׵/a;���}ɮ������bU?�Q\�����z�8�Z��S�w�@���a�D+x�nm����v��͜T�tva����?�2��L1��+pI�
�Z�m�k�����8]��8��1�G�aam§D���,�.N�夛d���$�Q�9ޏ=`<N2��or����7A�6�Z�+���sGF�����-��v�T1���8��RK��b��l_A�<b�[T�����O����2��p	��^:��)4Y��%E�zCmե~;��F^hND{8���ܴ��2�V�~z_���h�����$2�2;D!�ۈ~,��|UwX�Q��N�p��v��K�s�yv���z�L\�F�����"�Z�nm{�A#z��ۣ�=q�5�9��7�9;�.��y3DP�ԁ����	o@I��"3~������"m�Q�{3�!����_�J������H=i M���:�$�d�}��p~M�'�x�[��ɗ���f�|��F�qW]l�1Z�{:�����+3�+F���ux��7qu]_D0;�\��Z%���E�f�nS!��#�ˊI?Vj#��?V��u�����T�f�(~Q�� ��h�8��_��V�=�'i�u���Ε��G7!M��[B����23���|8Ё�u�@C<��76���x��o-AѶ��*i�$��.�1dN77��|6��Q����9���5�j��|
���L�2��D�n<���f������S�@�;D�a�?0k�W�9s�1�Ԕd����F*�Y�+�}�A]`l ZW�	�{pp~�0���`1����Њ\�/�D�*7QC��g�A��Y�q��7&���9^�b������:��,]��]ȼ��ͫh;>��H��3)OK5�����֓g �A�Y�C@ʅ�"&?ԧu�#;��W	�o� (�p��r�k��{�	س�pe_�����}1ڌ=$}���%���*X�ED)4��@�,0�$�F"��jx4�<�O$==+[����&����][�����Q@��T��|+01����wD3������\�̐D��;鳷������}���L���F^���<5�Wrt}�R7i��ɲO�5=Z��a&�:��x��l�->&2G���ƌ͡��v�Q��>u�5^A�w>����YWS�S"�r�ܫ3z�=�i`��}�~�<�]gk���".�Q�.��s��ːM������|�x.������$�K*��&��:Q�ad�P MF�Y�bm��%�I�a��%Y ����^L�:LkEa�w)�8HU����W����D�W��r�;�����D5"`���%#�4u�'	É�F��^_4E�S�6n��D�p��{����~���`�~|��p�<�B����!��4p^]y��d_����	�o6O��s�*���fR��V)�VF����c�b����j�í�w,X>p=3��͌�Q�oGk�|8<<y�y9���P�9Ws(Q�x���<�<����i�d���0�v������n�Mk���	O��ղb��9�o�`�-H��j�A�8���2��=��!�=��ʲ8C�(����O�B�PU��#�1��9\1ԣ�l�p�K��Z��]��Ȼ��M��j�F��X�qF�1J;��&>G��=��>f�!�@O���׌Y�i@�D�C)N[��<3�2������1�!����F����3�<��iHb�([-�E�k�gj�=i�?���%W<�խ��0p	�۾��Y/�C�8*�1����k��:1�D�&��� T�+��`S��.��[�{E'��K��4cЉ;��(%e��x�x����dt�־�g@v;ǭFF"���(�r�
��l9p.�n���(��lJ�B�oQ���geuoN\��Rz��)f�ˮTe�>�
(,���7��o���]͟���$�c�dT���.d�g�LZqեa���e9*i;�ZX8���I �hJ$؊Q�����N��D7�P+ȋTs�Y�4J�m�W��u�"��#��3�*�'P�)u���\z��O.�� ^����[Й�	*��}n	�;��޷��%��;�w�|���Ga��֘�픿�B���yak$M%��6|�>h����c�ϲ��N�����I!��l;>,����e��r�_c���0NM�E8}��9O*l?��_�M�7���5�b�Y-�<�t�u;I�0J|�!��[ә/�i�*I"�5�yf�����UFv<�{<A���1&vq��5Z �Sq1��K!����be�y�����"{�m��c��Wt�������?��	4�r<J�E�X[B�r�9l^�x��l�iپ到�l�m����i���9�l����J�,�h��7EDN�����bG���|�f���>�s :G�H?�Ĕ�l��I*}PU�)"�|�~Х�!8?({�/�4p���4��&=Ib�y4C�;b�$�#��NՕ��\�rH�\ ����v�1B��|܋�v��:�ߧ\����k p�I��⓹<�Y-%�w�w���3���Ŵ^x	��u3T���4�>�m�������fi���jKT���G��CA(�4(tܢ���ƒ��M���+����3kݴ!j��O��xM�_#�K�=��^�C�X�=]Cu�Iػ'/����:߲��F�6_H[A��vY�E#��
L=ә��1��X�cG!d���0y�Q�2a���=~ѧ�SgՅ�[\!)|��Ւ�\F�dSy���;]�uC�jv�������R+̏4i>w����M]���~��q��3�-2]Mʐnol8��sBj��p��JhBoC'�'z�H�ۂ��O���c`�>
2� dY�Ǖ[]��O*��kjk�������j�Q1�W���wG�$E�C8k)Aqn'��=>�x�n^�-NPC&���x�i�j�zD�(�&���������屋�>�J�Ơ��S�b�8/����0%�_W�R}e(�K�w�?�]Of��^ ӑ�x����k��u���G�(�oR��������w9A͕����7t�?��T�K/����Tj�p2����f��@!�q9ƉI����� �����j�$=1�%93��؝�Q��.o��j�!��7������0�����N������� �3�8M�����n��O2�E������;a��vC��N޽�qc�9�@m��� L,u:OY�}�I��*7)7����x�_Iw�RK��͌�����2P�����Z�6u[�l7n��R�(0�X��s�<�w	N�6&����B�Y�o].�}}4�o�b�`(�y�6j�}��^l9"ί��.H= 8И}�an�}P��ީ��7;��2�W��@����3��#(Cm��p�'�զ�0�V?J�1B�^�jS1���7$��>������Vgq��ty'�AJ�=������
-N������7�4M��G��X�m,�/��1��	��(?��:��<��qt�E'�7ek�q]a�Ej��`��	�=U� �i`<�i��{+�h�2v��5�|t��x�����>���t�T�	��\2Sx�j��k�xP"K���c�-�)�l�jsr�R� �]�E��I?��i3�k���bN!Q��L�@��s(v���^�K¤X  �:���1���s�k?&?v|r\_QA��|��}��'AG���K�|nY@�ܯ�|�tE�2CC7lV�-9d`���qb�z���m��V퀫~���I��lKy��ee-Ή�m�NktHr�h��*&q��JXH��MHH���h�*ǃu�������X���#���W� �㪵g��}��#\y�I.��Y�`��S��l='���<u��������>BY�ݤ�$Lmc�Y��<�`��y>QPa
D����E�i��0���siw��z��ܫ�ґ ��)B�3�-��t�.>?i�c��n��|���o�����{}Y[�)�d�7�k(X �YZ 	q��.Q���\cה(d�
�6	jl[�*��������?C�%���o�"M y���������.�B��?|e:���C�푕4�0!&��6��Ϋˀx�Y�<j��������� ��BԼrj�j�I"�+{�������3y㞬���x��<�RPn�\�:)���T�D�o�.���s.ʃ�E�p�+��*���[f����D�4���5y��0-V��I~y������Nkh_�2*��FT��Cqځ~�XLX2D��Z��Kz`@�7<�"uԇӆ�;,"S��~ivgh�$�tY���)�)ȎBH[ԇ
-�����V#*M�k`۝h�d�ɭ�Q�3������b�܈D�]Vu ��CS�a�0t�>T���n-h��fY�m��Vd�"ݩB��� S*{���̥������Q�T)�teAb`J��P���-�[,�TpB�%��ϭ�Dq� �՟�%��gQ��S��;'9��c_-#�rx���%A2��P�+��!��17��1Q5z�E�	Y[Sސ+h� EƉ����"��|�ٯ/��l�>e�1_]�l��LK���\�1�)ά�.b���.<�ʫ��ζ�)_i�]���O�r��^5��k2�bB`���V�:��2��%y�����\�b:��!a����T+U��؄��"��"���[	�q;֒w��7�4�u�k�f��#�����ے�Y)�]~�
��¥�?o�Q�a���5���M�T�l���I�]E۽�{p$��$�*���)��^�9	<�,Y��#M,���>x\w"�xڹ�����Q���q+M�E����#�g�k��ǳ�ƭ�¦ઔ;�:p�S�yH�Vj�����޼��6��p���"�2eI�O�
`�����ͺkvVs�y�:,��w�hˎ,h��2��@Ӷ �W�h�!�0_��9 ����ǜ:�k�y��s&g�8O+� V� ��� $���i[`������D�Ա�X�f�=����h��l%�_���.�{2���,'1���B�����
�7$����c��	jV�h�1��\}����^�tܔ֖9�G����]��g�%�hOVn�H����l+����/�p�Iu�v%'ԯbKU>���f�2h���g�a
�+�[�N�^$���Դ]���y��� O	��X��J(����Gװ�P�
�cR��N�{���_������9�vk]�2�?W�!�Z��>�v9x�Erf2*?<���yՏ_�W|T���k-�ݡe0Afa�pmDH��"fYo�����]�+l�b��i��a圕k��"D�xS��a3C�.����w�?'�jD�	3b:��)�z���)�I^]�3��H�T�@�"�g�R���m�3)�.�nf��w��i��2yȞ���UM�i~^���#/*�k^?��'���G�����=�z�J�׌Ƽ�8�b���Ϫ�-��EQ��e}��x�S1D#�x
��/�魽���ڳ#B��N�1�����^��ե�;_��~�tI3��w��$���[�ca[����]*���-�X����E2�o��6�)�@bV�Wi��Q)�e�Y	��6�})�bVK��[�q�j) ���=�1�q��8�)��2�(�69�^;/H�M?�M�E 6WF�{�tw�=Pe�I�ak�fcl�n$]��mY���t��\�5�	ÁZLB�Q���Cru!�1,q���v� �0�:ì�8̃���p$��m(�a?�b��������D�#POU��GU�kYg�`���l��cP}*�`��QI�Px��Z�U�^�;9��{,��+��m�N9���Z��ώ�KQ_�͟�v���M��g�U[�b���9�3��W�t���#�%��qV�9J�%9�i���8��"�6���4U�(`-��hc�w&�]�l#����m���]\�7�tF�"����������,��}M��+1�q 74z�[�Pl�E��7���[���П�K����$��PYh��6\.�����c�H���j��Da�]�*�л0�e|����� �c���T/҄���R��*�If�oi���Wy`r�t�v��OE˝�:��ƨ��4���/h0�`���p�iLP2���L�!��,;��A},Є���R`��X�l�װ��i��PD� �#|C[~{\��x�5"�'j���ϵ��M��j"0'��C<!������(Xyc����߻Z��+��M3�k�a�*y��8�me�a��bLX����D�ۿ��؅���5�.G�Ӻn��G��X=������>�-d��8� �y������E��r� J�NO�j<�Ç�z"�)��o�Pۦ��]���#{%�3Xb�%��y���W���קy�����"�YG�S0��|3���%�,`n�Გ���Tn*)j��p�g������8���U �͈GsЪ��b����W���,���\^ǶHXz��U<cN7�J���gZ;a)|�6��&�vw�p���ZO��J~��݂���%��k��,�YW?ϼ@iL
��������*��чtCW4�0�Z=�rԦ&k�5n����g������	���Y�y�F��V)�w�L�sߠ�g��GݔCw9B6���l�I��Qg����:�쫰e�y ��I�o�kH�;�{��x�bF�%�$�3��ھD��6}ۢ��y�K-���}���K�1�8r�b\���~�r����2�H�4�_�H�wի�C����0�m31�34AE����r�����U�X'\9����WY�I �����:R�4�4�a�e��]^0M�x��l��J>�n�*�!\a�	��p ýV�I�'��A��*����C,�*_�rѐ���ʄ��/|i���wh�м�eF�欎��^���z�	e�۔���~���	l��pRė���++X@Qra�����/�]�?u��q�(�!$�Cy�+�{갩B������0+��gb{�kJ&o#4��r��e����p;h�����=%�*����?T�:���7>9�[|�D��X9^��OP����O`����h�Sശ��2tl繎T���p��2jL�7L�S����]L#d�/9�*�{��"H�ex�����w��k��#��]�Q7=&;Ǚ|#�U�K��ex!w�k����o�͏�g�l������_~�a�S��=(�wo׳��._��^V�������8É���p�P��Qgz�Z����kjC���uS�'� �<�¬��)��|�e��Hٱ��� ��K{���xH5���a`��i�H�[KQ8S�� x�KT������0�ӏ>��PmG�v��^tqD�kk�R��Ӫ���;��ED>>���AB�Ҙ'D	��iB�vv��S�_%rc��D�����όV�B�U�/ww�/=>�Zm�c��KO,��`$�<Y��{��6��Q�@����e�#Q���.�\�˹>ß
����ĠQtr �}0Gʁ{^(��V�*�B7%sވ^��K��p�Q��9GwM�
�J�|G�H��H��,��d�T@�X���)��\����	�l+�z�����{�8����K�+�{�Dq�4k���P�a�Z�a~b>�ٕ�,��e�|�����l�@0��hZ9@Lߴ�]cc"�u@�l\/$�_�nJ,"%���Ri^�u\�q"���ٖۇ+�ܿ�0��Q�1����H�o��+D<�
*�;ށ���_Y��'�(��Z]���v��dC�#�i_�֟M����31~�(�ّg�ɫ*pr���iE�;�]��E���%� ��{g�
,ܡ�3�b��u��T��qPO&(��Oj�5��2�?,#`{��ۛ��d=�p a��sye�H{�"��h�*X�x��*U���ix��-�� $��>��>էj 0� ����c0�QFJw�:x���L��" f�l�C�N�+��o|�Ftk�o�00��d��AM������
|�,�U�g|�6�,�z�)e'_���Tqy"Q.X��!]�r�m��p}�l �+F
�ݗP�uP���Gw$�'o��D�,u.��kԤ�0%[l8�){���m�	���J_q���p��dѱ|�4ݬ���9�h.�r�H��J/�0��9��;�x^�`����_>\L=Dd�B��f�2�~��	�np�q^��d�hv�97O�Q^�g�O�' n�V�fb�����T)�Q���@=��Eҽtr�������V�b�õtS�
Kļ�s�� �Fs��K��+8Ѭ=\��.��3uv ��3*F�dI�PdP4k��|z��f��hgt_ڶ��m�X�I�[��w�c�J�+˥�xl[��HH��M_q�I�e�$��CIr,\�td��g�94I|%-�I�AJE��!�` ����q��`��&tq�K"p�R!�K)V�؆'D��We�_:4FvQe̦Ȕ���^C�����B�uW����N��E��WPi��ĞJ��H9�5.���ﲡ�_ /�V�"�:��J'��%�H�W]i�ꨴ(3��anB
yHj�:��w����Eu�6����μ�o��j0J>�FsGJ��zwb`����-�wА�&�/�Y,��_'q9�5-J��[�c-|[uI��=5|�I�}V�L]$ �,^x���4r/��65�7�&ߕF�%@c��=!�?���P�����tYŪ5�ߙk=��bCc�,*�j�l�ȝ�Y̑y�XPM=\����6{����;��& ��%Ŝ�MD�>Yv����\Z7|m!����td5(sn
߷o�y�*��wf����V�[n�m���$�y+�Y\����j$�?h�8�������#� �ԐJ��w�o�O*�����1���;�i�GEs?�(9h'r�oH�
Q/z��Z����e�,���x��2u9�Ϫ��R��j�;��
�@�����\�L��7VS{��H`�]�k���ȍ������P~B6}��5%�,������;�z��N�O�EW��*	d��tCa(\s�O)/��h�=s�<Q�{����v�9o~0�s�ډT3�����y#�1{�d�����������&�&�`�6Q[>��,�� ��6j���H�R.����㋾�7"`s����6�F2H�_P>�����#��ۤK��r5���}}�sP6܊��֑0�qs��/G�ՄFNvΨ�57��l�V��^���Y[N�P�:��4t��韻�{Bo�ߗ��E͕�X�\�Z�9���Iu��HgB���ǐ��V���-�Z����TW:�'�b��� s�q�k/��Y�����D��zY�-dk�x@�kiM���թ��D�aH۔��KGV���_�x�����V?@�k�V o0�+p�? �?����e!�ɿx���;�.$��AHK5�8P=��)�~Skė�X�)[f`w�X��;A%��=�����SY���+�W�5��6og?�	��*�H:�H�̉Q��b���,t�$�YU��]��陾�A�v.����q޻��C޹A��k!#����BM�.�v#Bd���Ӥ���F`Ԫ��{"�ξЀ*�����T5tX����� �A����f'��E�A
-�_�����j"�a8����(q� �ﳖ��9@�=��	����U�/��]G�s���]y��ϼʟ��U��V�j��QI�fw��P������B�12�~��4��:�y����X�#
�r�:]vK'2���Zz�
6����$+W\�Jt�d[cI�i�xl��
D��q[#����J�Cu2� *��Ү�D�}7 ӓ�'���~�Y����6��k��GM��m���њwvX��8�B�׹��`����c��c�C��ha��I�"�}��v��of1��ڞn�^�>�ķ�����ܶo(�1l�O�,@?��֚l˰*c�����
�c9�N�&P �7��=����X�#��9��KӾ��3�fC����k�����E����=8��-@&^$�	��F��.�lq�l�7�o�=�FHnwz� B�h��#��b�T�>*��IW^�ƃ�;l|��W�A�=k%��3���ꑁ\xm�St�"#U�)E�+ƻ��,I2����Iޛ��9��,�1�S��������]��3e�'�(d�TR���w�u�27��3�d�"X���[��Z0�_�DOHm�5\�άg��R2�X�l$X7��
�,��[���+���-��L'fJp��3,���䉋�,�fΖ[���>��Mv_5A.Cs����ٍ�ss��>�+��|^��@cg\�%T	E@ i�P��l��LaKafG���\��EȩFLd)Z��qZ�o�^ں`���0�df��8�z6�0g+�	��"�D�� �Հ˨�Ţ��]�)�7y�dvR$�ޓ�ju����D�S�\�<��δh3�w��ܙ�3q��ɪ�%�a}���/ �p�$P\��t��G&e
�u�o����f6SS.�k���s�&^�&��I�V�J��z"��	b����8�sxl��E���L�8i�Z�M���Ok����d��X:��QO��V@��}�T�ŃI�FJu+9w:ˊ�M{�7�r7Uu�-Hz���!a���0�a*�wee�bu���9�뚼^�V���m?N�/�NF��n�:(�OG�>����xd�H�h��BBjs�|��'ۯ���\��I����X���
�т�1�BiG�q�2s/�q�.Õ֗���`~���`	���N�
�ŻR�j��ſ��e���rxH�J/��� '���)E.�qḁ����1	�H���
�����}��1�zP���=]���itα��ˎvX@�����g��Z�����r�$�����"��J_����7�!ձ��j����SM�1����Z��mM����x�e+�U�"�翪�yݬ2
�
�Ǐ��"��u[��#+���Qm�sF8�W����S1�S�j[��sAx�iR��Ȼ�0g�&��F�rZ�&��]�@yج�pju�W8����Y����͝�D�|�s0|�ا>��H�V<b:�-�8"��>E7OE=U�z)�n�v�:�0�ϻ$�m�mV-�$�>��z�L����<`�
C/���,\F
��b�k��E�������&�~g�Vo#Ӯ7��N�<���L��Q��zQ\��������`U���?���A�7����L�OkE*�2.s���%8@��oX��".]h���1�p��N7Q|���-�=�[����OҐ�PYٰ�Ӷ$�=�C����xy���-�w�m�ё�"*�I|�!�'PlUD�r��G7�(H�$���4��ď�Q4��0Qn�F�B��Ct@1��9�f�a�u��,(�
�C.#j�̸Qԭ��y�Q�GA�QT��mf�"��^*d=�Ɂu��:Ò�B=j��M��KUGd�Z*����iτO�����#��5����?��'�7���I�EH�ʉ�DP9[s{%%�� (�[�/��1���pb��Dr`�Q+&�0V }�=����tԙ� ���¨�#��v�^�E�)Iw��&}��|�T�x�Jʤڼi�Mބ`o�l[F+����$���y��V{��M�Gӓ�!4��
/��UE%Qc��=��b���}�g�
QK�`6�4p`��q��b}�q��E"�Y�����ȵ8G'�~�9��1:_Y��[��,�j�~���e�;�!��1fe�e@Ĭ��@s��a&W���7������+tGI���HT����QG�!��O;�քO��Q���J�m0�;\d:����T�C�����S�����ZJ�qm���������{ry`o�f��E���1��̳|+�e����ڋq���5�3��������N�|H�}j\�U*l�t�S�欌�ܭ���3!��I]���8�&���-��2[:nqJ'�r��ˡ�V�W�$��I{3	S�1�;!���>�*�q6Dv�ri�����Jl,P�ȹ���n}Fۨ�.�q�X��'35�D;�T�T�Y���'��8��ٿ�ߟ|��_�BwN�e�==�ke��5����h/�Lһ�er5]�X���Nz\��߉4z���#���c���<��О��	�r�Ա��$���&����$�kF�I�Q3�f�x�%r6)�gB�Z̄��e�0��Gq�6�-�0
�j��D�f�>��VZ#�j��{z�x�Q��~���;����?��jva���'.�8�킨���� �Y(K�Nh&�N�y�>U�s��xS�>����OD�r�|@�E�ۡ n�0�,6G⑫��g0��3�y�2ȇ-��FU�s�FH�s��}i�rb=?�Fk'��jeC��-��Q;mO�@�m�m�w>2�K̏UHk�������ѸɖBX����.����r�ݯ�~7޸oN�l:�����0Ơ�8�ZCX|�|�4ve���Y<�!0��� �&�ً�EvrC'�Zb˪��ȍ��:>b��eĴ_bX�/�n��y�I�]8Ֆ�5�3�"F<��_�$}���+�C`.z�G�1��c�f^������㕗-rZ�P�p�v�췅Z��V�(�*R�㝡gq�4���"r,��������Nۣd�&���OA����-	�������[m����E��'��h@���?X=�f^12y�������K�R�
C�!5��<덺�D��It�;E�A��Zs�ARt�69�@�5�K`�Pܛo��`t���+�Pt��>����,p�s�Ů���~�(�8��Rݝ�qH�O���\~�*J�;FM瞙�������4}=DXr�`�-4`��#���0���i��	NID��H�Yf}�9�Ao��g�|�f�9�XK31�{}�㉚�t�C�����K'�p-	3g=,Oɦw�u��3KD^�B�gXƗ@ߘ�ͳ�)�9I�4�+YF�Q,�G��i��H7�A���O�v9F�'g����_M�3ZtC��]�SU0�Y���/%q?���GK����~�Tx�A6��Q�+Ri7��I�$j�M,�|w�@ڲ��^�@���U|2֨@�D���� "����2��%b4`��NG%��F/��M<'60�9���$�3yI�qZ��$�h�!�ð�74Ә͆�Օ\�ۯ��H<���ao?��&�:�Xh4�,0`�]o�A����<u�+��Bw��&�K}��;��ة�oꨫ�S��S����Atm��z��}�,vF#y1^2l����F�[��n3�[⻈9��Q7���E��#1E��FT��v�#[p�t_��[6� ������@A�����x��I����]L�f��E6�K���I�Qn�-OW�����
�f��4� �t��rpA�)�^:OU��zDD
��n�;��S1�iH�2;~����6�X�xu|�L)��I��DN�t�����u��e��$�;�8�g��Sf���m�cggC�]$���D�(B�t�ä! �(9�g�p_�e�a�	.(%m�1�1AV|�?�*�!�?�&V�o/-�����j1�yi�^�m|��z�
1�����!k~��W`�pn���튜v[�8�s���X�FG���ŭo�$/Z��ɆW�&��C�q��]�,�.:?ʣN!P,Fn;��k�-Q�@o��Э(�\��q�ȦR��vg�tʒK
�K��";	�V9�L����>?rN�
��}��1Xժ6/i�)���7h����¥sw��գ��hTm���s"B�`������	Au� �<7�N��B`��'��������	i�e�/��d�q�	� ����p������;����*��pq�;щ=㰀����wZd�������@��\�1�1�S�R[<6 g/�,�m�:"Y�H]-j*�N�c��yOȗa����P:#���&�N�Q��0�TiF+J��a�0~�O����Mݤ��)��D��(�/Q*QZ��:̙���=���ܫ�k@v��` +��%#1�+�wƲ�e�gd��$ �iR	#�����T��$����̱�°;�s��ڎ#���ֿ}�B����F�R�l4��[���]�'Fh��,&#�k�g���\>��o����y�
vrB��5���QG'�L���V��v�Ɲy�I۠�7%=�@�|y{�Q�3���ǎH[�x�psŧ��
"w��08OLfq˧5� ИF�tT"0&�xyb�"n����7c1�r:|����_��^���+K�%d���T��I��ދ"Q�kЍ�2��	��`���F���Fg��p@��C�7ɜG�E�+��ޞ0d�$_�!<S/����׬�s�8yoMWN�A���;"�h�����E����]�{���Y�Ԉ�^��^jL�Χ��c�k�~�*ޖq3����/#º�cBQϞ�� �Kե�$��U>I�����,<�Wz���;Ab."U��f*��i��]0�B�����H�g/'����|��|�r19"�e'AH�"��;M+�0⎀�WB�wG��,� \�#Җ�"�RPQm.[ӹem�F��#(��H����
�����~
��]j�𰙏�'��-�cO�V���`�g:���gWA�qև��մ�I�1A�n�:�1Hx�
�vI֡�}|�~!�vT�Do�h4A���A��ed�	9D�upj=uR�ݵ��A���Z[�A'lQHO6$�$��9�B���"=E'�.�݊Av�.���"7Alp:G�~�q�g�$Ǌ�h�hb�$����"��&�y�-/�^2�KCCIk�f�D�|/6޶sL�܂���HkKD��STz{0ѯr�0��>�wщk���ŧ��z�V��$��l�3UʛP�����rʻ�������[o�Ģ�tZ���*��q�A��/��r�1]a�Xxy�	�o=p�T�>T&�gKe�Ps
�H��G�\��Ҙ5�[^���q�
�[F�v�vX澾�p����n|�X	E\�q�5h�|铸4��!{t�9�i�@J{U#�F�֕j����	��o���N�W?��J��H��CL�d"
�[\��	`�ȋ�eM�=nF�Sqһp^)�"�N�ϫ�xlGG}1@��x��Ku���&=Jz�mE���]yL�����(�Ǡ�D=d�S�M���r˗(oN���@�����;j�8B�;H�ޜ�zkX'��R�L���1T�>��B9k������=۩J$\t��O� ��M�ˡǢ�
g��g��ļU5��t����O �����B{3F6U�;�]	o�e�{�+��X}�1����UsU�~���n��#*��!=��|���l~������������q��@���<�7��kn�à'ڸ����c���2��"f���D���&�Xr�+��&�T�x"�|K�}%����S��O�D�J�V�4:mͨbp�G��0�P��PAf{ �tg/ǀ+ �S�0hM��-���z�pO��,�x�/"Z.�Q�{�����
��y�[�ǲ�WÓ�͹m���s���8�T�r�}��-oJ�tC�3}���H����0�����)B��H�&���/��8t��2aTG �T�@_���G��y��r5`)_FN	(����$
�H�d	�G6a\;��ϻ#wS0�7��8tt�q{�" >���"
t{�;�gd��������uȕ)1A�XD��ݏ.523{�Pڕ�_�Csc~0XLh�tb�^88���'�MN���� �5���]�����!r��	���܃U�,�_;��0�(ՀkC�����s�c���sAuG���&G8��`M����
��k��HQ���0�����s�8o�D�J����t��Y��',�"��C���Əiz�E${�r K�д&���pJ�?�Cl��!>1�M��I]�r`���P�CT��/�n�Ꮲ��X����*��v�T3D)G�0�Ð�n?�+��u��{�hw ����-Z��̪�dy�b4 �����!���?%\l2��*�}MY��'�J��_вW�YQ}���B�Ȗ��̫�0���U�Y3��t�HI^(�0>>F��s�����;<���^+�$l1$��T�I�^!�;n���8>S�;^?�GC@��Fm��wlQ =���Ƒ��{�g�:������T�dK�����-��\%�I\8T���}�q^E��7����3������=HV�>g[m�,c���ع��{l}OgP����]xF�`d.f�1�U9N<1$I}v��܅e���Pͪ�=��O�'��_�u�
�~���[p(}9zT�r�т�W\�r�'��6�J�Ŵd^�����38TW���	�?[�}���lX�;�#�\��u����r�)�d���j>�����DO�jC��+���f �e�}�)�Q��m�`$+���B.p��~�Q��
�j���B�o� cs����u��Qq����)d�M� �?��CT͚������*'%���vA��~\���>ћ��iF:�Ռ�X�&�`�ڌ4W$q��|�.5��(�Y� +��fOxtZ�-��Ѐ�u����<��$�}�b�!��(A�Jk ���A��r��R͂�|��ѥ���˙�p$hYT�ɟ`}��ư�K4ד�r!�弣_r�m�Ek~{w��k]�>E�Ͷ������U�wt�L��N%�|(�����ǼJ4밢�g��Sɞ�:ȹ�1�hm���X����-���a��NSi-��!�ӧ�Fy�SDW4���±����6~Y}&	?'1(b⚻1��Ӳsܝ�eK݌|ܪo�幐T_;�\�B�w�u����'B������gs�[ �6�O9�xDh��?��a�V���(ft�7�|�H�U���W��*�%C��Q��1��Y֞%��3��h����^_� :�o^-^�1����A�M�K쿔{%���k|O]�H�V��9�a��(�j&�4�ƛ�f�j��)�WI����m�hn���;��n��5>�:`��~f��lNT6�Xbo�GʳG3V�6�k�E��a��X��5��:�(��5AH�AKP)$��?���Dx��I8IJ��zk�t]!bf� 2������a��^��������~=/�2���&r�$�����c�ԃ_��+�u�hO �	?�E���C�^{�)�<���C&I7S�Y֚|�ΈXY�Q�Pu��f���0�nxu���S𤢾��:s`/5s�?V�ŕ�
�M6Cv�~~��BT�5J�Xg,�������"���=�q^��?�QwS(u͈jkܐ��o(&�g�dn��l�f��u�c��z萑�,�u�����a�
�s9`��܍�>�˝&��}9�C�y�v��TAK^%��\c��7^����\�pr,*k�(�L]I1��vϻ��3�F[	������o�UC�/3�up�Qk�^+ws�܎��z�r�Ew�K��+)=��W�&��y1@ؖՖU��l���jX����u����_"b�'��tXw>{�z��;\Ӓ�����U`:KQ~EVь��� ����)�8�7g�-����&! 4w@l��T���/��`��v��"�dl��X��Ī�����y�6���SK|HH���t|m�9� ����
�DKN��4�<,�
�c����)D��k��*/�,k���7����K�O�N��֮�ͣ��q@���$,e��|7��B��[R��P(�������"����+jz�Ф'jDQyibH�x(]���� ����߃�D푍�)���6�~�����d`�������H���n��Դ�7��\��ZT:'̓��� ����M�9�9r��-�3�۫;A��{�χ�vZ��z��)R�<�+e�/�ԩ����#�G'7��#muE~|�SiEڿb̜�m (̰���ζM��bD◵9�%X%���<JA�Z���mMl�@i2���o��Q�b+��[~����%��,���)kP(��/��`����`��*�K�X�3�[�3�JҤ�Oej�������/�{?rM3J��94���$������n�ɫ99b��{��P!�gڽ��e�J�k5�c���mJ�7���ɟ/N�����\�G�d�
�'��!�b6ٷh���4�/^�Mj�Y���&w24ӱl~�y�\�\�P��3�����҅NIdE�!�-
��P?y�j�D��a��p|�'���=C��p1�$wLbK� 3�˯�O����󈈅Ri�� ނzAzb��G^1�z�0�CY�|���ZSמ�t��xi�A;�"�җ�<g�y ��mN)EB��I��kA�O�#ۢX�o�-e�vl�ݝ@7=a(z:��~!H*�p3>�I���O���݁���B����p�[��a��}�q���>��]'�{���&�f��-j�m�͘��a��ѣu[#��B	�b�q�r��g��V;��p�4U��`"����`S6ﺽaM�Gm�"ԯ��Ő��3�v�o2�X�0!Ԉ�&�� ���FI�4���"��'�|�uԆ������w?���*�T�<p�c�\L��;[��%kQV�U5z4E���`]����(��[�1^�:��ݮ�3���u�.�lS��o������`9�4���ieN��j�Ф�3J`� v�4���+���*��ER�[�y-���l��`D:!E/�o���#;5���nu=�z!?}*%r�}%�,d�σ��sx�|v�{j�6��g���дܧPH��l˄%,�D�����#�;SL��`]]T���AF��e50	��^z����P�_gkjrPCO_���?��˯�|q� ڋ��l�q�ΐ��U��YpȦ*\gX�z����s?��D[Z��d{Uy��K�}m\�3���=��_b�� ����5��S��y�?�I���������R4&��=�.�K��Mt��I��\T����uVT�ތ��U�N�q���5짞s^vH�$���\pL����I��z&��S�,I��d�퐈���<0?�W�9wp�
7��탄�(X���=~���ه��"�N��%��2�&7��Ӂ�	�����H�p�ˇ��܉�験�i���4PLU�[&Q��j(hxne���r)��5���
D ]yD-�,)�`�N���� |k�4�����/n,=���BY@��X�����#b>8��U~�Ԇ=ӪQ��͐�AVU �Β��	,��p�k3�����z:���(����e�X�p3�:c�>���]��2�V9�n���P�Wkm�VB�10c�k�k<��X�47>��*� +-�=?'��Iwi��}z'B�5P}i���m�|X�E���ğX�f:7�Q2^ў��¿h�_P����'�0��.�Q_ 3�)�`�պ+���&�K��2�3v�s�Knw��e��kz�E�#��Ƣ���D��P�Fd�.j'�6�>�@���؇��6��z1��x_� �Mؗ�}��l~�7R���j��w��04�\\�A���������!���uDDt`�n�KL��%WF}~�ݙ�p �*��fw%9�����Bu�u;��-�k?p�v�m��>�������s��i�Q(�+Q.J��1�%�u.��,-V:�@��)�Bv�/��mG�����h�U|;�,u�m5�M�n'�Q%�k�X�_6h���&���>���1��D�ǝ�zQ|h�)	s&�Ր��56����:��'�Q����6m��S$�
��hnR萦鴿�����Kq��~�Y;"T�qp�x~i�?Ze�P���<� ޛ��/�哙��̀�e@ԧ9Fm��HL�_'Q	�9@[T`(�Ч
M	j�M��dL��A{�0����R��O+��C�g�ѷ�f;�ݲ�f���E�T !�婝�&6$����
5׭:�n�:ǲ]k��|�����cy����*�zq..9������i�ch��H�\DF`CO�J��xs-�12�.������\6QBRQr����=�.�tܻ��`0�쁟d������G?������3�߃�ɽN�2�d`6B�d�C�Q�m^񦔍UY�1���NHco|vxhP��y�H�~o�Y:�ؠ�0aGI76O����T���	�PA�u��hx�M|� 6�V�olP��-��!Z��i{B]'\�S������_�<�I�,P��'�?�#��m`�]0�A�':��4#�<_~)+RC��!WP�.��V�A�i�ծF����D�sM���|�K#i�|آ4�����&�:M}r���r؞
G��އ�����饡�{<5�P�s���rVJ;IF��={���u��5�}�k(t����g��[�"���'�~��eY#ǩ���6Gg)i��|^��VQ�.�}�h�f��m��c� �f�>{��4��F�
Cm������z\���DA�J����kG���f8
V�K������^b>�����m:�����R��s���ߘ��B��HX��Q��=�$���Xc���:�iO
��~�OK��Ҫn��ZO��J��)��Q%�S\C�����Q�M>H��ѰaC�l���q����y���9��Zo��U��6[��Q���Bg�DWސ�Ӟ�]&7b�jO�
>���~��v
`"<��9E=5Q��,_=�� .�'�����M�����|��G^�N+E���S.X�!3���@�9\�N0���4�I������/���	1�yW�glռ��2��͠�SK���Џ�VO�-�	�S��'E�nj�T\���G��e�M㖓wK�*;�K� �sa�p1l�o� ��ڞ���`i-��jZs��]UO��E(l�2T������BXj���Tת��9��lPA�C;��8Q����f
%��{f48��u��/�eH�"�Ȇ���d��/�R�%q
�C�S�6�z�����v����7o~5S3����g��i����G�:XC,���l�H����$�	oB�H�-��*`��rݜ�VG��Vg�1�u��[BN�5�X�ܶP]c�������h�@w?�ќy(rd<�SF��`�NF1�K��PP<U]��$b���/��3ɠ�cW��� :ȣ� M�����z�/�7��+n�/�����s�A �c
��r;.稅7��������!$�(X/]�"	ӹ��$qD+���2"?w�H�P�?���`��������C������J����k�%A���&_[�4V*�mYiQc�ÛY��B�[�\uZ��Z�<s����E4F�F��]ݽ������p�ѻ���#8�{9����� ��Y̩����'ej���ۛ
B�Ϯ�m��ڽg��Z�_��h!(�S�?�t��u�̒S~�fM�:��UpY���Y�����dW�3#���}�uػ2Z>�0Ͳ�cf��_%'�������O���҇�s��1�Y)F)�`	�P�ޢ�6��5���c��&w��٧9!b���mM�f�܃#������؈�Ng������Q*\��	��ͭҰ�X`t�6���DH�<Q��O�~�,��g�]Q��Y��+;�����˽�b3�d�6�N�Hͽ��Ґ��д�}?T�&L�=��8��.?����]rє���5�C+�n�ƎK
����ٷv6����t��d���
b}�v�7�9���֚s���Ӽ��jB͓k
�.m ٌC�����k�x]B�f��Ex���&G�w��Jz�P�,��G�P,ȝd�����đ��>����Q��~��0�N�W�|���VH��\.�SBF�Z�p��eO����=>�K+[p�*G0�ѿT`
$ʅ2���g�E[81�p�d��Ղ��fgt��:�2�Q���J�<���X��s��Və�d?�a��Q� �ܾ_��"�����f�sr>;�nJxEV��±��m��7"B�}@�{9t�=���I�j�l�l��10?M��{�E3As��)ǽ��ý����\�0���mJ� &m�qU�Q�1|J�J�>91k1�i-���.���	�K_u�"�'��lP�aPZ��ɚ�[���k�(�m7g �D��U�T�,� N�y륋0�U�N�gzeS�q�2<H��@�k�증*�e
�_	��U��F3>Χ��d �~��.�R1'C� ��=�)b샮	{U����P~��2%�L�cv��=Q��ߎ�@dL	�+	���ߤ$&
r��3��/ѝy�LG+��"�< ���#��|4�p�s��.��ڤ����fD+����A�����<ҟ{EԶp4zT�1^�ލ�#{tϘq6�i���yY?�Ɍ6!l�%�Y�@�܀�[��X@�%3Ao�W!h�4� b�֎�4�c�'���h䀦d��9��}ĩ�0�O�j��������ҕ�� �}߂�G8d!K%��3�2V��D1�:�xl����C"8!���B���0a��!Jr�o�s6J��2�!j���N�����K��2O�����cԾ���R�����r�Z���a�_p?��lF,'��k~�s�d3�z@��P��qcM��e��+8�9E��j��ktq��JEW����{^w���}��pb����r	�9u�*��+L�,9�:��}��0�EuM��[�����R膊��P��������G��=x���f/��$��>6���Cȕ�p"��Jgd�@*Ň���hX;�Y�Z ��#�Y����'8��&��R'uM �72%/��y9-�����p`�e�s(��U��Y��MzJ�PV�Ŕ�NW��a�y;$dx1�˗�5�����)Ŵ�虻-�QDu���&�&�e��yN���z�>Ƭc�L��_�
 ꢪ�\��^Շ؇LK��M-��q$��>C5��(""U~Lq��Q9�gG[W����~ ��곞�}��1,�;!��w��}�L̚K���]�9�
��|�_l֜=F�W�ժ�kkmlӞ���ܝ���.�_Tx���ym��G��HT��'�L3[���y+m��-�2�u:�-�B�zU�&#� ��?�AP3D���# ���ٍ�4C �/�NRM�rs��^M��|�\)=����^�g��t����J��FV@�c#Ģ2��r7��������� O8��/)����X���*�f�W���D[�����x_�V(�tU15�MV��{��~CZ��'�;���Q)ב,=+���#<�\�d �}���a1��@�z7&m���U�~��4�ڨҿA^i�Z��%�3;�][Fw���E���C�Ȓr�v�6��9�{��V}�S*������W3�fq	q|�x\Oy��L�����Q�i!tJ��{B�&�J�-��B?�eG���ާF��R����' b��4V)`��~�:6�x'T��^W�9u�tɑ|0;Q�k7�:Ϩ�	af6w�m.��ե�t���F��C ���^nsQ���6�A��cq�/\oU<.mn[gI�Oc�oo��sw�鯫e�Hw�e�����0Y���!LOI�BAC���y��&�j��9A�I	�)JI�-�����έ3��W�i/�3������.y	��My��3։.��6��@mƵ�4���[���\+��9�P		Nf��s���B(��ް�-�FV�W�`�wU�p|�rpfV7R.���"{����&�Am 2#��ä�z�Q$wi�3�)^-p8�f�KO��<��-��_��~�8\^0���d9P�߅m����k��<1Y ���N�w��1A��>g������		>��0n)�
��zI�Q@��sT.z��[i���b�~�S@������h��5�@JmQ)M,iŘ�tB.6/wBC����K����)I8zª؂��i�AgQ@��Jϋ�w".�#9�l�"%�Q,��N=Px�LL�� z��c�A�_�%�)?����[���V"�G`RU����ևKG/ͦp���nY"9���0��D�3�Kk'-�$w^1s�żE�
)����%�9 3nhZ�����8��J�LY����A$`+�&��PY�������0?F��S�\�sm䠝$�le}_QK��E40�܅N�1��}D���� �!�.Q��.�o��&E�VK�s�|Ww��)Gd�l�'I%�]+_�!�~ئU�dK��0k��5s��-�i���52�MZS�s�����R!t��JԢ���Y{`��I�|��6��y�ӎ�v�&'ʛ�Vb
�E�;Hy�,�+������L���tj
�����9d���d7���ZT���G����s�E����x�%��,S<�_��ȉ��ub�Oa8+�3R�q�W��Cs�f�6��W��)�)C��7
�W\��2�>���)��l�`%T�l�ȑ�s��3Vc�У�U�Þ2��xrS1�3��p}}�EX� ů��-X��OR|G��N_&Be��ý�ψPRldV6�_*�+��k�lNV��p�<��_d�	Wʲ�U4�eki����L�M(�x}��eC�]q����GXB^��TwW{�N �@�S��ߗ"<`����;X�+6�9���@'�woN�hN��n��'X�lB?k;��<����ظ�9���˰��,?:�Y�6�n� >�	w��{�5g*ʶ�;:e�UQjd�6�x
�B���7S��o�<r�!�#p����ܶu����c��,ؠ���qr�@�Ì�A%I�5�ម��k�do�sI7�2����8;yht9�f��w��7y��3���R�p�}��z¥�O	�,�mH��g8}w��i's�|TD1rL�옵��Q���X+$o��2��) �摒\���	Ä���$T���
�m�T5Vڵ��yJ擃���GZU2���8�<yczݸ�6⌐cf�Il�����z)�S&�$Ψnj��~m��І�y{c��}~o4�΂b-Ř�y�ʮ2�@���%��@C� �Ѡ�\[	lx��4q��v�^T���<(��
X�3x1 �
y���l�����|d�P�Uy#DĿ��&�3�����t��d�ƢpaW�1��9�2�u7vY���tn�&��`[��,a��Fn	�J{�������u�蠙��-�+�� ���B0a-C�f�P҉hЖT�k�Vg�[f�����i��,���~_Q.u!�>���u&]����R���g5�H��R"�.���Oa�}�iF�V�sl�j����O�K�p/2^�j�`3�buG7 �U���İ�\�v�$�������%{�TT?"��צf���)�a5).��E��R%Z�,nN�Y�Zm���h_�/*)2V��-Q++jw-���[K�;���A5�<_ �3'l��I��b�m9�Ob�� �0�?�	k�M�N�������,<%���Y�a�FȽJz�d
����:ڤr^&\g/K[�ޔ�oRq�>��e�$�06��6�0M��͞�sW���6`���a�>5'�(�>; ��G��M�8���5����#nIS�7C9���3AcE] &�8_=�񿱽o�K�)�R� �/����e�h� � �*�nS�@��?��ó�@<0ª ��7��6����H��������pv�w/<�be/>$<o�����A��i�D;�󏅙��Pwc/D�/���R��I ��� ��l��t�}���vz��_+t)�T�,
K��m~M+{���#3@xe%����
;oNN�:�B�����1�sW�US���ڴ�B�+���i�J�~�}[� hG���U'�86�[*�i��j�ɡ1J��ji�lf+p�G��II��g(OEURo�OC�p��m`ȴ��k�	�BҍH�� ٛ䏶�V�po�R��R�9"e�"`�﷉��V�ve�<b��z�Wo��;�5����5��Ԏ,�� c�
T��,��(��Ģf�.E3�sV�XL��&q��ŭ���es:�
�Rxel���:��Fl����`�4���+t�$���嚇���^2�xRF���I��;�~1���H6dmP"h��*����w��uD�������NC[�sb*��g�o����Ԝ��4��3���:�>�,ٙ��â̜ςWf�%J�f�0����9u�+�B]8�� �|���!p�����0U����Qyn!��}V��!�:�B����f�B����G����1�S�����U�^d�ȋ�0g^t�0���A�艃��m0��
���Z�Q@�Gss�^l��*7�N�ȵ�X��&$ι�/L����.[�B��n��O�����>��J���㙃�82������&E�<y���#���#X�M��.�����;�U\*����I�0�<&X�TW��(���{T��t%��6_��$K_�2��7f�X0&Rc>�S0�Z�}KtH���;O��U�c(���i�؁�1Nl�J-�+,��&R·ZQՑ��8��E���jԀ���i��PS�9��7�HǌC���Dk�b����o � ʚB)�eL	� G�g�St{o��)Վ�j@��4���y�$�F��̽c���� 㰐���`R�I�������2��+�-�yX~���R������Q�	字G�����h`G^���������k樦Q�j[�H	����.� ��%Bp7�Jy"��@V�%d��d�pi̤��X7����p3��� ��"�^�U��<>�)>���������*g�tJ�hI���V�Gy�}-��ƫo�T]�<}��2N�wL�<���0��S̭LJ�+�d~�ۮ�q\zMc��]���.¥�q�(�cQ�\;hh�}�K%�L��x4��&,�>��_	`a����b��5��^a�F"qs��~̠׮�C�����M�!\0j�aa��K��<�g�/��P���d�_��S��C�F�bs9�}���4�Tܫ�"kdj�!^�Uձ��5�L��_IЮX���L��g$��\�u��ӶG-z�ȁկ���r4�}��LA-�3���q��Y�?�aPN͢�l�|�<�H���?h���u����z���;��Ta��vU:���(��=4��M2��QN� ���S�p�P5���\m-v��K�}T���i�&��Q.{�YH����9��3����hH�n��t�}�V��ͳ:$q+�#M� l�0IT�#=�F�{B�vt�c����S���v`n�P���;~4v�c�X�����Uɽc��;�;�W�C��V�K����/�n{�H7v3�\W��4�C�-dG����3x2�Ɇ�UY��� .�,}o�p����!/U?�&��5�f�������vJA��&��ͧ:-�{Z4eq��×~Nv���QH��D��=r���/��	������<���>�:��.�H�s��cNDZH%LW��Гt58�J��n�	�8���;�a�&��z@JÃ����ണ�ҴE���х�.���sx����^T�9W�!��z>B ���̃��1(~����5bV\��"~��'��+:�)Vu�"#�&���Bg���Mg�Ǹ�1��q7���U����2##���l#�<��%{�A�������=Z��K�� )a�è���#�R��R77�u�� $�=�F�re��5�|)Y0�?Ne�sc��:B��*҅	(�SFW�u�E\5#�&|9~�-�g^I�D��\��u8���A�Ѵ^�e�Q�r����so���>ܘ�E캇�_�����&-l�NG����5YE��]s$G��{9�o�����-[5�@�A�&~�.�w�<�X�N���d,�<���9����g��\&B�O4���<�PN��q�D���"�#C���Gr�lT����|�gE*[-�����"S �I�	㘏�Ǵ7{�2�^(��ȇ��7��J�"�xJ,CDZU3��Q,��ʞ�P�I�J�L��r�P��)�s%n����5YD���Lo��n�%V�A� ���G�
s�J'{T>��1��E�c���x�,qh���o~��w&��2A�P~�(�����&���5���hM�6�/�9���#���S٠S,y�9S+��Ԇ~O#]A�m����_�uՍV��/1׭���-�q��+������~�:=�ܚ�kq�ϱdh��(�=��Iy��4�a����Z���츧2��*HE᭄U톆ww
����]�[��ؗ��<��߾�I���& A��A�,+{x�K>��	��7��#H���$ԕ^t�M���c�):e�b�M����T�̣�&L#!���IŬF^x��p���z��!��,xF�
k�6Q�$�=�u���O��ʈs}�HO@`PdN�rIA�Wo�0��z�M��.��׉����.��~���x�;�U�,�۞Ą���:T~,���H�Ȗ2�6��|�+���d�����{w�P�qt �؝[�TP��vj7�βS �G��{r�(5'�|��/j�DᏕH�w�JG	��.�����|߭7>�Q��?�R┦"aI/��|��!�z�oೡ_#	^�& ��4�^�.�º�<=x��Gq�y0�@*(Mz�<�� đ��2�����̹���OC���)�%���b���B�lи :$��qi�c��=<Z��Bb!v�X����&�$.�&;9��&�z^4��{��\K$e	�sŚ,\�aEgq���^�
�]%Z?g�[��h��P�t�Ԍ_�&Ǖ8] _ ŬX��.�۹Zʖ����D�`A^�t�x���#A�r��s��qw�\j �0�v^_�5M.��ϗi#|?p#���\�8f%�K��_R\S�tx��2�5��v=5�*��`� .̼H�J2�2p�	��t��9�	x��{	�n;w��VT|؉3�VG�Y6��'%�	�)��-��6a<�{��gvv$G9Nzf�\y��@V�����������^�W2��D��-C�Ũ`�"� a=`�LՐQ�읹�(4R�Κ�B�L���KAo261�.n"��Ə����cM͍����,޲ll�\�hn����R�$يo��A�g���z�J�g'G�� �Ck1BG����MF0��d��ƚ��[�8q�糜��~���I��e���,�����E��;��OP��tECz�/�,��X�|�j�Jjnj��)zh�+2�5Z�r��z�� ������X�_sq��_�C��.�B��JTA�*��m���l��@�vL�UJ��T��x^J/G�Ձ(�� �ԣ
�����f/�~0�s7m<����̠�����:��xV%
�,�iH~���-?���d�W����Ɓ#�vՋC�L�W�T�#Q�+�!�/SZ���T�Fh:�yE�cC~ܤ�z/�&��fn,�w�o�͛����0ps6�l����>�]��}S�-qrf�<�cv���fe�;v2:I�>P�b[�We���=V\[�z4,9N�"�� sW����-X�U�F���HJ"��XNl�'��.'~i8��W��k�9�������Vb ,�K����kۂ���N�&�;��y8���&�4Ru���p��2]��f�:�؆2�z|�H�C�jv3�Ө�~�S6��Ǯ��i�}��7r+�^�e���h�a�u���	͞��y�И��.+�T��%��*�W����x���{�n6����P��;M��N�N���Q��,�_@�FÂ�t-�8d�7�I�A���[����:�V���X������W��L�$�\��T��XѺݠ�:�}�� &{J.xB�-����Kp�*s��잕��kF�^�V�\L޶f!��Y��W����N�N�$7�Fщ/)�!��Щ�zT��o�[�t���f�,B��´� ($����g���9�|�l��-"�
��X��`������ �3�;�`�0w%���#�E]����F�T����������8��x6����i�ؗY~�h�5�8���<�����0%�m��/�W��g���>U7���d���65D�J�Y������ǿf��ؙU�lLC�8�� �D�j��Xb�p�Oʕ䉧��0O�W�.Z#l�
�Jl�ݤm@�-����<x2�&@�9ӭ�{I��hVf}���N!-��ޢ���o�f�aO>��`n�haF7`!Nq]�dHTB���S�: ���oL�њ�#J�$*��@��x�kՊ�]���ʁLV�?̹���O��l�?�ʳ�z~�P�Ӫ����@�Q����i�������'��}@u�� �^��<�f��V�S���9�T��W��̰U��,����c4�ou����G�;
Y���TV;�)N�>[�-�Msr�X��f��'��Z��h����&��?�ƯN�&8����@�8��������Z�*є#��~��Xߝ߭V�{ݥ�CN@�z�ꐦ��E�T�-ӂ�*��"Ru�$����s�xKg�!a�|�R�.����u:�j]B�!b��?��(�[�	��6LF��Ĳ��.
���Vv���������;�U�_Q�pZ���d�ǲ�^�~Y )5�_�p��f&�j�i��e���꿱���A�8�^h�J�����5��㟐�I ��ك��$v���	���s."h�Q�5j���U��7�C�Rv)*�w��'��8:�3�aJ3=�����XO$fV����P�� ����{��1,k�lG�2�U(�pɭ}	6��7PcGv�e���n�*?���Ϫ@r�~p̣��k�^�N���bB�Y~��-���n�]4E`"�M�̦8_k���'J8��T}��nT�+ϒ+�ׅ>��]�{lo���W�����"�����-�dN�Y�|�~l��B��Ӡ�_�A	1���N}�����(�X��@!���m���y�m�1��RU���7�Y�B]��R<�t.&|s���<S�>h�k?,V8a�j�Rw�!�g��_R g�c�2�NRN��[�Q�#�!֎��[�6H9�$�u�0�6���x0$øJ����T�����&�7B��05pRH`l"�\���Ko�\xz �$@-1*3y���j�˓�ir��A�!/! �?af�!�@�b�ٽ��u�d��lb��[b���o�,��`�Dl��Wg�P~����f�I`�qXȺoY�"i�Π�Y.A�@t�^4ƘS����Hn=pS`�_K���e�8m��s*5W>��}}H�������Wx����o4�ҷ�=�Z�}�9��=b��ׯ)FJ+���fB˵�Y�s�ЉuF��*@PD1oH��\�)�����wh�Єp1�K��pdmw���V+|:i���KmQ�y�ז���1F=���#t}���l���4^k�y	溥�4O�b4*Qk��M��tx��:��m]�U�=�Ms�3�h%X�Ɂ}]w�9 V։(㦥q�އ��y5B2�J��(��x�K�+Y����@\>�c����'D�f���Ӳj*��t�]��:�}�e��;�,��D$�=ۘ��� .���m�v�6�Ԏތ(8���T0����Vs�@����Q�4�>w�K�h�AO/��a�OG���*�G��5
��ԥ��eAcTQ��x�Ӂ�F��"����JAV*9O�;6�l��n�.{گږ-�{;  'A�W��,���Od͡�bU�1T�L?t)X=�O��M�HnnFLuEt���'jD_K/�m�h���w�P͗I%�[�L:���� wG���B�b���Dâ(O�:ڻ��x|�>˜Z���!�+^DY�ѣ�H"|�4pO������9��qg'�7��*��U�{��(�_���#�b��A�����M��S�}�� �?Os��dA	��zP� ����ɶ�)�'���af[]\6���ￃY`� X|�C�MJ�*#�5�-�\��?Vw�+WLq������!h�N�C��/�'�U�A]�|��	s��ju+��u��;�L�a��(�c�d��G�$���;0F��kY��Y�B�t�)� %������g,O1�����_�?eh����ܐz�7��_�d�u�Ũ׆�2(�omEd��q�S��ɹЃܗ�5P��F���`>��k_�m��M����J� ��gl�TC�*����"���D�{_��u�Oπ��;��o�Rx���oL"���\�>mZ+8 ���0��7X�R'%��si�96�l ���XRĔ��_�<��w(�HƊ�s/�v~����;P�u��2�4���kQ]� r���	6E��ִ��Xz��k�QX5�N�w��!URD��_p^85I�qw��eMt��Z���-�c�<K|�2�vB�V��É����Y�
U?@�v� y|Q@��ѱ!R�����шB�����(��+��>�TF	D�+�h@K]����t
�o�n��!���^�5T��M�++��U<L#D���i�=7�T�1�9���x�TRG|��gi���G��@`2�\(�+ PT�`+}%=�w���˅����G��W��o��U�=�U�T���
p =�p:Q)�8{W*g�q�/jv��/��zO �;�����
������Ig�0�]�Μ e��̑�Z�kW����(�����KM���|���PJ��1�`0�'.�uO����b�)��i|u$:�u��9m�@�FV�6��xҭTg�@��k� �?F^�gG�A�P
�
G�d�ܧ��!u�~CÈ��C1�zѿ!��\q6����=J�{�w�S�xn��9�xb��>C�"�3Rj����>��q���_��è�Kt�����8��_ghT��n�<b���E��_g%�/AƊ��q7]��AF��CI�G�Rh^�.�D#|ĕ�Gf�JF�H��w~w�'Q��e�Ke�`ه�Q�ߵ�X���i���.������<�Q���h��H)^��B� �5��o8���ޏi-��f�ծ�
��^��f��>Y��S��3"�+���]�v%mЧE�Βɤ���ڷ�t�
b�5� ��*yj��L�c���n����D�+UG�C%'f0j��������e��;ό���]��:
L����4Wm��ߩ��!�NBi��]��z�,���~���d�B &�.p' 6L2Lr"�����V4��'���q˘XQ��®�E/[�/v�,�����#:~y��Ȥ��C��$����Q����W��xN�m�Gv�ũ�@��E�p0�H�Cc�aKFb�h�%sΝW/ͺ�cB)ռ.�.��h�j7�������7=���C.��x�~�[�(5�BJ����V��5�	�e��$,����U恿}3$P��˻it�ě�7��:�eZ�c)4 "���n�<UI�����h��d+_�i�	&�5ۏr�4�ӌF�	�#½��;2U�r�`F���/x��=�)�N�qv�H��cP�=��([�߷��8��>): fV��i�}���ڬ��X������l�
�zB�A��J�3���ۈ�;�?�@�rv � d.J����M���,�
�0�8�m]s�|���������;��4�14�k�N�d|��8sR�#���/-�-!��0�گ�)��������sڻB�i`3�r;�ʏ��ۃQ-����>��P��枣�����H���E���i΁S���,4Og���ҧ�?��wwy�)x�Tur��ۘ�~�]�a+	D��O���@P6�|L+�үf��֠� ?��ΌQrQB%�om!+�9h���|�m<.���#��u�32]�x�Mx�����HZ\�����jp4P�t�+uT��r���ٶ*���l��	�&����PA4=���y)�J�����T*Y���)a����G��J:C�͛�'���g������)�X��,�5O�*���5l�ǂ�����Љ�nt��a�s���&�5�^H�C�V��>��\���3��͍ǉ}�DPr�hފ8:�4�]��݉="(x{ddAd�6�\W;華 >X[�zZe���N,;�4���[�s-4;���2�D<��$��.u ߛ�Ԕ HP��c�w8>H�	:� %���$>�N47��C��&��K��Ф��p4I��H��H d��p-��A�ѝ9a�g�����u��0F�<�mr��*��'�Q�����{w2+����/^�١Ƒ�9M'(J�	�&��;jpA��|B�}��ϡ�^9���S�5lӹ��n@�N
���b���?F��
�4�
J��CyL��v��Đ�g�c�p�&�������`̻���9���N3/���:�9N�{|���Փ�1#�íT�$�5d���m���h��w���O��b@)�ZM���5u0�N��D$��:u��i�B�N���!��@��ėEk)Fw���Y2���j;���aUvO8�N�#�Ց�o��9�r�=�����MN�6F&�>)Yhl�5���I���� mm�ޔ���{�r�ݸf>[���.>0A�*uZ�[��=V��%���pW�)L6a@\�h�1?�*��Ó�C�q{Vڪ�&�o9�(�'������W ��I
�M�)�[�s��u��a!�z!g|�>!��X�_�Q�2ʫ��A{��O��g8Q�R����F��!=�Y:v�$.�����= p�N��}��ո$��5�$����_oe�ʕ��Z4���#"�u�N���u����d��0hW�U�j�=&iY�����  ���I�!EkZ��&+�y�+|�Ld~o��J�f^5�����M�xI�8C�QqAI��7�j̸Z��Z�kÒN��-�f�u�a�C1��~D������,���
J�Y?��t�+4<	{����e����{����0��U�V�p��d��V��`�|�7�S�T�+t;�;�۞䰩C��i��K��o���C���;�_-Fv!�h�4&�״�!�z��1��]�! h�Ɣxr�{�64��ġ���J�VW[�h]����bLrN�uk�p�cr�5\W$^6�t���\�-�,lX��|�f���kc4.�Re�l���jO���f�$�'����OM�6�!~	>b���fU��df����$�"Q�J�	��/��ɌK��-l������uh���]RO�΁B��Z�>H�����q�I�U��Xm@�{�Ρ�m��Ӱ��l���9���}B�-�5g�̘3��s (�2��,�%)�&B�^�X%2h.�ag�+n�#����,3e�}�`�6�u3�y�vLk�c�H������8��=�
բ��c��jC(���n,��f8.�-��XP:��/�)|T�.;5�j>�}Rf_%d�<����r�V�G��$A��I�}74�[���7�C�c���+�J[��D3����Ccm��j��9�%H�Q�g�4Xf1{PJ�;����1��\y��Ŕ�����J�&I��P�$	K���{������>�-q6r�8��t"p!��&P��^N'JBC��g|�Lx���&���W/�rn��w��n�W���P�-J�֯� ��4�at:̛�邖QO�.���蔆F�<���k�<K�eVSWY�6aU}��[�Hp/���ir5 yP\6����|#�N��;�szܭ&?`aSI�`p����j���\�e�>�d�P��x�)�:��z�TLT
+#m�����&۴I��Ma�:</��_�Ն�]S��Y��
����V:�����[b���Q���$�N�葤����S/Ӱ7[��fA d�	e-�|�M&Yp5� ���)!3_}Q��A��7-=ӽ;)�@���+��	��7�&�[����5���ͺY���y�%k�?�U�oue�59��V��:b����:Ț����_�- "�׺"]`��A��I��e�Ttd�J[ΪZ����3^�7nW<}���U�C��C��y�K�G�3�o�w�x��2Jr�j�&���{g�t��S�N1j~�أ�(Zfݳ��=���G��L�0�+�B��tQ�虌�F��t����D<���ã4�wm���}�[��A;��{�+Ɗ�Y�|Ghn��n^�Q�9m�yL\L�����#U�����4��I|�y������P��j�z�Oiu�n>�՟@�Ç�S��2��8���������Ġ�#�b�\і�����9�"��V'��\�t����'��6���J�>��4t	J8EF�J���6��:�O(O�n(m�yA	��gU�fP�YZ=c��z��mV��^ɝ���^�z�ҝsڳ��]�5�9MS>�Q��Р��q��LN��J���_��Z�N!p)K�4D�	8FGY���9�'(Oc���Fϋb�mQV��T�0)
��&�^�!d��]���t�K�&i��wc.; ���d7���/��\�A�s'�4�~uGbg���� ��.��x|7=��{w |Ѵ�P+��r�D����<���n>��7�詢Ҏ�=�
N+�*�=U��tٌ���;�KM�>Y�w�.և��J��h��Z��#,��=��fM��ת�ڤD����#0 t�!���|<T@=���6v�Q��i�{P>9�Wn�԰Z)ܘ�`Cڛ�w���ԕ��� ��p�H(JB�e�x�ғ�\�K����C��i͍����1��	!j����A��
u�f�ٝ�c}�ű�dd��C���4)˕�UN�]'����c�II~�[h�	ۼ�/#"�Q��!��K*	�E5e,�(�/1�Ƞ%MJ��sp�<|7�޽Ҩ_$���9����jq�ǋ4P�ʍ�j�0>�uhy���^��_�w�󳲨����a�<���!�k�X�3OB�>{Y���O�+�*����j8y�N�V�:0u2(����}[�EmEd`����'K���������6c ��(˭�*��h[{�~�ytzvW�]�I����[0�a��:Q�Z�S�����t����j���8���z>Y㖧lƓv
W��J�T��y��Sذ�|2�!=��������
E�Q�sI���D��澾ʠO�
��{�N��vp��?�uS�j�F$�o�9�<Ir��C���&"�c�pO[g=�O���Fо5^Q&�9���T�L8I/ն><%�H�Qf?�#���<
(��M����EG�b��M]�h�bE����׻./��P=w�=���:��Ԁ$4�S[�\<�	��ɖC���,/_��\��:%�e6	�aVrƼ�%��+O5K�3dV�����u�hZ���׷�y�3M�f�r����7J�o�w.�~��6e햣��ӥhr��J#���P�#~���D��C�ۙ�k�g��͟!^��qoO(��Or_!a�xjT�PO��,�'�|�[�d;W1l�?T���9� ���K�}ȺwN��yg~��Qq%���R�,n�R]�?(h	��Fk�A!GtA��	A
�@�c8��f��s�ܡ ��&��^���|J&51�U�D	�=�^ ����I��b�l�g��*�b+f��3*A,���K�t�I��0ȃ%Ю��#/�].�8&N��C�QI���;^-`@e���U��GL��Z�U�!�h�������[��+ѾZ����_�������B�DhK[��T3% /�p��n�n����%Gx/�"l�o�<�!,!���D�0�.�9Htzs(A��)��we����0�ᯆ �RK`�$�U��ؐ�ʗO/'Cs�$~1�$8��x(R�>#���C?��\I�0�c'��-Ό�]�k�ӿ�N/�u�"��՗��b��=g��T;F��h3lͤ�(����aOC1��Xl���T퐺1�e`Ϭ\�d�:��ji�F@ʐ���Jg �c�&��@��8���J�]S\�|��o�.�AD���ba�#����X���W�����C��!j���Jʡ�hJx���#9,K�������XN!�W�0] bd�R�[
<�<���A�8c
�Klߊu�릗ɣ�ǩ`�����!S2��U���,'aw��j4�,���q}Ґ���nb�:�ȲyG�����Wv�&Ad��5p1�kƴ@��j�[0�МB'�8}]�y�'z��R"Ut�؁�,�#�04G���hIT�y-�!A(�L�GS�dF���l��W�3�@�MQ�D�$'JxqR'�E���e\� ��t��A�>tn���:7/�=�N44�]滂~5F��`�7?�5-P/^���k*_���`K�s�*Ǖn����A��(�����?Y�{@d���8AY���4���\�8,J �����F(h�c�N��}��J�Z���S���inyAD6S.@�A��>����:�D']��2`K��Pf=��)�%�������V����~$B�=-f{���T�������ݡgĹ��W]ӹH
�<Y��k:�;W,�+�)�}��������o��L�M�W}�z�Y4t�wd N*�	����(VJ�["��ZrM�.Q��N��w#��f�qՕ\��(Q��|�g�/1�b�M����N��y�υ�e`SWJVP��3 N�� A�X���=�z%�T˧�6H���j�C���*�^�K8�3È��	�}��!byX�4��i�տ���V���Y9�мg�sZ���U受xӹ-��&�ݒJIaZ%^��3����Qξ�O��[�s��gj�I�h�������s��7�7+&G��~��]R��I��^�^ @C���Ea3/u\��N`>"8ɐ�$��֪�W[= �D��  F�B,���4k���ZB��n(K�ǂ,İ &��N��"��7��н���h.��T�ʓw`~�)n�J�(�t��C��BC��p����L���a���?�A���89	1�
��2(����g�gz2��щgC�@�VPSS*���[��[��o.�}��qץ�z.��X@`k-kֵ�r�
�,��16dNX� 熝~}M���f�~�=q�]8>�>�+c�rj!��;E�,�,�z�2�Ɔ�r/�%�چu�S��#��n�
��:&a�=���WFe��M	���ؼsP8�YS����1�9M�|S9)�9r��$:lM�6���s��g�~��S@J��� g�7�����Q��q���*Ź��ygU��j�!:X	����Rx=��ޓ:H??�UQ0�4�}�5��4k���n�)(u�?(�x��6K���%�	$���q�鰑.��A�J9�O�bZ��}�A3��6���9��G�sa���r���LDD��w�;b]�Qإ~������ud�o��y���;�vbepW0�=��ܲUH0�����qru��ڄ��=�=��'��*6^<,���>�?�O^-j!�m��0�C0�?<mSC_���ףF�+�'��	�4�rU3�MYJ����a�,����<b��c�0��K��TC��s�%��a0�+��|H��@��Yє�G��9\::L� A�uɒ-����Q��P�0�2jN��N�����p��;!���{�v�6�g�0�,?8�޹xW��ڐ����C������Yt_�R�uY�ѱ:r;U+��n���zE�+Ϭ��J��,5V"���	GtK ��ڃ���G��܀���k�����:G��S�>�UL���)��;�b�ٴh
eBM$!�E�t/�� 1��l����@��e#��Qsإ%82QB�*�T�<H�S怛9i�{�>��vג�UI��� �ױJI�A�"F���J��`#�n�)�����y�+��
3S�.�l��sƾ�;K��)Ss���}�_$С�q{Ic�=4\	u�n����z[�z ����+c*���n+���ڂ�,*Q��㰢�@FH�o�1�S����&����px�NP�- 4	�X�*�CLx$�:w�OU����!�qٓ��%�=�Y.1s0�Ԧ�b�\ߠb�~�R&�K�ߠ�w�GSXp�ޱ���sF���������*=P�l�2*��K�'�f�#��j�ڒT�-���0l<|����H���0t #�B�L|��Yí2�
25C�����Nr54��2S)�:>�&��2�� ��;�y�(@���3|�Hu1���&!z��w��JB9��Lae�
2�m�a�S0 ��Q@^��L����K�<��\�»	���]�4=�׍�$�G�ȭ�}~5��a��Y2^�����8�I��X���V��L�!/S_�t�1�o61pN�X��[���7�h�V�X�K
�7
D��t�����H#1��a��lp�)�y�%1ƨ\b-lȮu��Rũ5�z�r_�~hUz���Q�%cy��0�=9<x2񶎜 �Y��Ii�J�t�6����m�&�����ܧd}:j���z1޷0m
�q_�.q[5̯ y�>�4C4��RY�θd�|[�
�#�̣�"l��Z�-�R�KT�"�`�`*�^ ���bH������k2����R1������=�a*��2��$�����IWc�˃�d�4|�]%Y������Ra><x�,y���Ȯ��:�hM��$�/\�
���I���um^�Z�����/	�1	'�X�]=�I�fmo
)S�������%E���V��/��\;Yfz�w�<���,�n؞�D���jT��٣�T8
T�X�Y��#��s1�0w7�(G
ok��Υ�
|K&(,���*ZmD3��;AN��<�k�Z����@�)C��j�6nY��B3���ܡ��ȆO;Q���)��sz-Ӹ���)N"�O]�'�Km�1�f=&"�m�]�$��@���%������r�Vq<�B�q	��\�LKP����g���$m'��0�V�Q�7%�QZʔ�ٟ:��W�vޝ��[���Qt�'�.5�z��`�֖����^��\��?ܬN����}/�?�͊N�j)	���2j}�4Ņt���@tc9���˖�1�;�Eu��p3����/DGt/k�#�˨���M�(.��a���A��T.T�}��p����f؇t(�@k���y��;z��=	���@ק��t�p>����K�ɕ��E	O�Hq��O�$�������q��ʿ;z��Cㆯ��ϒ�띪�7�ʊ�P�aD�U��)���ϻ
$�G�?jV9�-V sB�::�s�H�nWC�{�j"nǇQݯ��^X�8܊���`fw��<��&��ܯ;�kz�G6�AQNƙp�����;e�<}�j&ۿ���v���]
Fw�C�R�g#��G z�r��ū�=�)��������9}�_�t�}��:�0�Y�����X�xdCW�  �]䮶M���t�/
��RV�3�/ �9���L[Lfu/�#(�O����g���̯�D	��^�^�ʰ�����OU���;(��������1�ŭ��A h�t[�D���i*���6�5hE���c�UN�r̤_�V��)��q���I�<�JY���N�.�U��m�2�,����;�N wE5��90>C�?Z4�(�I��:���jf��R��T<I�e����fF��\6z��ĵ����i՛��J&��;��a��V����8�Ʃpp��%יр�AU�������̠U�=r��
i)3�����\��I.��=k~j��D_�O���JSnʎ��{g��y�����2!�������s��\b%��R���h�R�0H'��Ci!�ϻ���b=	�WyWI֦ّ[�����C2��+V�+[�:�:n&P���'���F��U��>� J+.Ԝ5��ؗ(賻������~Q�B�N�}E(=�h,��e]�xWksZD� Q���.�Č<δ="*�H|K�"_���`�ѵQS�b��� ��Ap.A�#+ޓ�9BwT19�6]�0P�!��(:�F	-����>h2�G�?���Ln�W4M��,�r�J��K��Z�PdȀ�J�il��O��Yc
����B��ÑN���>m(��wv]�Z� d���O)��3�C!�����n*��QW����z��t��:�v�b��S<A�*�W*������]��z�2Cx��pcRw�����d~��B� -�l�1�_m?z��;�i�Y�6���Z���╝���>y�]#��倵3̍�� �� SP��x�([�.�D(w�d�<o]��ԃ�Qi#ϛv�]�8w�gw���]��?\m[�������,�q#��'3����b��p陯��kCGR���C������HKΈ���u���Ɔ���D��x��"��9�3�4��6ѱD�QwC��h�\|A����Z��h����=f��l�支>X+�i�A^S]�f�x�1�8�$t�V<�	������J3�ᐐ@�Iù#O�\����M�=�6�≱�Y��'��??��{�W۬k�K69�٨��P�8�ר5ե�ۖ�\|��/�[
 ��^�5y��F��0��2E�g<�@8:�؝'��nʵ�vM��V�I9p[jwQ�B�._��)��4��+�T�`�/gE���H�(9~ �gk��i��'R-��lS�7�W���l����/�~GΙZ�k;ChM�P ��"`�i�*�[�� �Ľ�06�6h] �l�0���>�u	k�׈vY.�,�.]�7���RbmV��/�ǹ�L�ϐZz^� ֑c�Fsէ+����zHM*�	��e{()o����.a�u��v_�Ё�6~BSք�D�c;��N���Q�o<��9�o��7a<�E�"�` ��q�n�,Ht��!�I��� ejD�^1�^2=q1����E0T���h�f�i�+g�U,%Xe���p	�e��1,����6�����v*�q�3�y��v��7̫�P,��G��NA�+�lR�y,�{�]w�������?oA�ɎړlZrU��`�K��g��i��;GЖ�G
k�4���#����j)�D�#��tM��*�ѧ����#o[T���i�%B_j�������.9����L��;�63�֮S`F�5��+�W���:YE��m`��:`�qw�2���h?f����	�d�����f�-��;Е!�l+���1�),�N����g�H�W��1%�"b�x~ɚ Z,�_X$���ȗ��)�[}�B�n�U��nAqR8[3ƨU���B�m`,��[���9�6�~ǻ`�*�y��� \�:�>/	�V��e��/h4O����^!S9�~����u�, -`��M�����X:�C�?}�gOW�G]b#��Q�]�X�C�Ju���P���o@´�@"�z{� ��Z��0��9�Wc����XvH�]��*ª\�o�F<_�c�\_��4��{e(�� �0����"���RQ��SR	~���.b �!�'a(r��VǨ�d����%���jNh!8�n9^�$N��o����ʅR�*f�Ĥ^�|U��w�m$R�葏Eu0>�	����[��ѷV���96�
֗��\8"o,S���ѧ�o���`,D�'�"���(Y/-��f�-����}���,�����]�|ү�s�|��wK&�@tfP�������|hPN�&h8�� [�<�|.�ӷ_�f����_L"�-4��Qj�!�+Hw��\�����-#zo�6��+���澋Z�%ˤ��^�o�� �4O��K��,ґ�I��5�m��=VS�̫�U/�m��Q�@�q�^x��+�vLy�;���-Z g���\��-]���
�:�@B��Ts����0c���4*�5���(`�Z۟���������&�SQ�v���f��ll�7Y�
�Ѣü��h)?�K{+aǯ"5^y��U�H����=����zH%�6k9+t���3���=-� dmo��Ι��	�e�xa\�c�mLa�"F��C�6� c��5bԸS����B�+��I���d��CE��������&"���DwN5X�D0�Ӗ4�rc�mlcKk�7��� ���3^>�Z�T�چ^�=s�c���؉�2xp}�b`�P��2)��ԁ���L�y?��a���r��{X�s��r~�7<�	��� v�WƱo��3�!	ZQ��nyq!gh!��"��t�H���f{�,�\q>�����L��lB�3��@��Wn�r�����<�0}���'�0g-��.�=hȒ��+��"����B�O`B˓�E�5�xR��tV�+��5��g?������7���Ȝ�w2�2#Z6��d����SQ��O��V�E��@��b�P�Q��V�q���X4�$�.-�ԌY��{�w�Bl7=ѼE�f[ZU�Ϟ-�hS!+ .��zI�ם��ьc����"�bs�,r&f=��;��t�
7)N��ϛx�MrQၦ�Iz�̬�9���ԭ<��t���3ꐉ��6f�䰕�;��*y��q���?��#m�>�%�Bڽ�YA8��|}fb�N¥4H�uqb�k�h�?,�foŏJ���B�ł�CX�`�]�<Jߡ�o'�7��;���`���>�����ē2�چJ!�ė�f���e�S� �L�E�ŝm|8a^;�M�Ȣ5����>&�3+�Xq���?��X&�/�����5�/��}o�l���s� d���ϙ+�_&|�B�{�:�����4G�Aٺ��[�������^�g� �J�{�3�������WE&6/KC&��H;���.~�7N�q뿂;Og����Ki�餙� ����	�I&�ŞL������c�:I	� ٶTښ��ZЄ�6���G5�s�܊2�bR��9
���1�߄΂i��^�>:m>��Mr���Z��HlA����ʶq��K)���л_#_�%/�侐ou�n��y{77
��֞C��4x��S��SK�J�}$� ]2�0�q�Y��.S9��Ws�K���Ű�f��"��0
�Ǟk1i��ZJ1�F3��(�N�gג���0�M����yMJ{�w7���:;���A\�� FaG��`�.����8��D��]�' %���'ź{��KQ����g?w�;,D��t�c}7��Ĭ1���Q��-�p�4����#D��j�ȍܞ(E�]���^��lIm_A�9[�jƿ"��|H�ͳ֙�55\��IY�ο��ʿ.��*������_�?U�ѓksiS��5�Z�nR�$P�20z�c��m6�$���㹎7s��0�7Ǳ������^��f��З`��}���.�<��^	Ŧv8ɱ0:'LX���]#��P��EQ�����&u�:���z+��x �����m�S�����{i�WWR�N�PgfM?�����F��E@߯t�B�eP^2S�8(��UoQ+�\B!X�!I�-��%��@*̂� ��X.��x�+@�b���d%~�"h�0Z���bp��c�!�n�ᒞ?�/�Fl�s\ey�,j�!:*���������a�$q��LA���YS8dL&>��h�����t�s^m@�-��1�2�� f�������A϶���V��զ?]��;c�EKi��G���	�u�k�A�^�.o����	:�qȑe���mO����{b�"=��t3�9���C}��ױB��Je�a�5�V�߲�3-��=�����z[�E��{��#P�7�! ����0\A�Q���S{��h���!�XjJ�l��{������_LP��kW"��ձ�O �9�&T�X�X�{2GF"�3���mV~R�Z\�xj%����WA�y�lA�;��ȭ����橙�.C�b[�<��W��*�v͆�3"�~ek��4��ĶY�m�
K�ʹ5�P���i�%���e�5����Q�O��}cծ4�
S��9�E�\�e�Q�H`#�^�)6r�{�(h��噧��!gh^� �ܘJ*Z�E�֢�2������n�ώۏ�<q<�����ӷ����1���0`iϖ&'�RqR�T�!NTVY���"ñ�u�,�Ȑ�?,��mz��$Z׼��q.�K}�6��9I����6�r_ĉ*1��P��0��Z~\L�c����hГ�䗅A��P�W�N]ޝ欠S�I�"����������?ՉBdpl����k9VAK��q��Z���S����g�߅e�������{#D�,�2�;X��A�
��� ��z���`���F�a���>r|���\�m���7x�OB��`��-�o���������.�8 6�g����ތ~��m����M���Gx�U��}(߃��`1Q�k�֓����`p�����x���&��tk�|���v�e�D[<ᩌ���K2\
���,2��sõ5��_�'��eM r'��R� � s���GQ$�4}!����Jm�?�CH[N�SPZg/��3%���ş�(����+$�b+��s/b	#��<��Υ��(j;�5%'����Һ���[��z''��L��q��0�x����L�1$�zȦU�38��f��s�ji[��D�w�Ҁ�1�E|�Z)�X���&���2Gt��2��f}�� Ԓ
W�DB�B�%���(3{s�^{�[�y�Ь*�e�����_t+>��T6�=8�e�A�g1�'ީ9BU�:��N��J�[�d�&�Y�,,��R���<��u�!��B/�,|=�d �Ih�;Ưj� Բ�M3蒝����d��\�!h��L���4o83#�Q�}o"�Hq�l�B�9 )I=�*�<!���!m�vGS�L��b�lǥvW�rMI�w��J��!Y��p[�`i]�*��m�K�P���횙�)8*r�FD�P���u��wn��m�1���r~Z3W�h"��欐2,��)� ���(Jx������̗��7��)��s�q�sl�׼@�臵�~�->Y��-�lTe!�ܙ��rmEc:�����meϻ�L�o�[�8��1A1�d��((:&M�4T;+mp&��l�	���^[-�Δv샘��Y>~i �J���Vv֎��=��%z�i)@���_V?�e�&���������'iRi������·d��m`h�%s���e
jHX��E^Ā�V����w��}î��>�A� ���`�W��YD����!����(ysIF��g:R^=h�5�g�k��ŋ��G�|��+M/�BT�6N�c³!L��=O�јuSo�֣��®�-]�6=0�Z���U��g=&}�l�!]����i�;`{���g��P���aQ=����v�9�վ��2{-׿��I��~�?�Y�ғ;)�nQ�3���yNRUQ���p_w���d�5���`E`��n�X��`��Eh�-=Y�K�o��♣F�����,~r?�ZBL�Pz� ɏ��Yy��\�����g��D����<��o����]:Œ���N���&Y��#<G1��Cڞ_��s���+���>Ԯ�E}ҁյ�m��R�fy��X����r;IH�x�`ʘV �J�j���m�%��z�GRz-��R�Π�u���_�qy�Dk�PHʴ�:�H<��Y!~T�,�	O��ݷ;�<����(���8~�`���uKԝ�0����o�: YR(��Kd�  D������<���N�BgH¾�C%�$�r�l!����L�Ǔ�=iuҹ0^�O�G7�f��R`���"`����Y"�e��d�$C�J�;���j�{dJ��G�Wj)@�)��|����]"�-�f�A7�Q��a�w�S�f��7#�L��"��`�9�~���#Nv�E�O��:cK�����������=�n�`�]p���A�s9J����C�q��1��}��\�͠_��\�R ��@�ayLY��]�M��j�Z%Z�0"��𧣺��bLIq�؝U�"�.����G�i8�)~q��>oG�����2��@v�,u^4잰�>`�[����,ƞ��(�p�6t��oe�2Y�� /���;r�^xGz�l���*@=z���!�x��s���^c��F����n�7�v������ k��@P�,��yk���o�>�t��N���m<���?��]6SqM�u*�C�e��f�ӠU���ӵ�z��#h4ӷګj�<�Uv�:fI,
E4{�*8F�͘�Y�#n*|M��f>~��`p�<�G�wa���-�2@��V�3�t��9vZZ��$��O2T�9%��y��;{���JQ��r����w����i����uˤ"o(��ʤ��*i]!�|z��	1��1a��Έ�փD��vMf�X����0��ਭC��Ƃ�ݧ���n�����\��Nx����8�{��W5�q���rBDp����+�Z�u}Z�����CX�1%�y1��5g����w�2�$�W+�T�[�cd5�*��W�V�T�ӝ/ha,�x?��\/��tUr���PH\nb�׌T��
�]Zyy)���c�';����{P��rZ˼+�^�x�����&$�)V�9֦�=i�8���^�r�׹��4m���`�Z���.(���,-�١�b`?��@��Cg<����fy���y
�
[��L�֣n���q6��=�_���
A�3~�=ŵ�'�!1���jm;����x���U)����Q#ǆ��Z|���τ�."]��"���0�4�r5%I�+4 G~ஓ���n5B�͌��:#}Z��^�w=Qzż�LZ=�{� �<�af��œ�r��m >ʽE�'����@1���k�;Щ��JS�'U�#'Pb��Ll���E��Ƈ/�� ��#���H�B�ֳg��5?��x-�D��&�۝�?`CU��>)Ꞃ��E�����q��\}��O�X�Q�~�|I�"p�\%�	 �b��..��sص�ध�7���&>�7Xg|�N��,G�Z�E����*"�T�}R�=�oM��z(J�t��A��5�;�,+���Ŧ�qF�<�����?<��+�����@s�͟O6�$m���S}����F�����̪�?˥��P�e����Q;�wV�!4����ӆ�e,%���@E�S�Ĝ+w��_���4������2��:�K�jIn�frw՝�<P�0+��tĝ4���B��	�,E�f8E��k�/wL'��\ð��KD�93���`W��b1�`lw�6�/��a3\�l������Gg�	!1��f�iy�U�����"7v�l�IĽ��p�b�.=a�U�Je�����D�6\��irq������Ԋ�#a.%��,t��:����aiڬ�q��,u�����6GKi��y-?q�����yK��5[�,XL-��H�m�W>=��qØT�5���Z�T�q6���`d̂z�n?��O����x�N�@!�%r,mI�}�W��n�����Ξ!=��,������|�Yf��ѻbnAW?
&���*b���F"����Lr?��H�]�Ր�5�W��O�y��f޿
NM�G�L&uĸ|�4ץu�]o�����ʦtK!�ȡ��PuH��G^�0=~xF8�4�ʂ�+��b]��\��7�z�*�+8���4<y�c�߆'��O펍Ė��0r+�S��v�l��M��N꿼���,GI�ɮyH�$�ZQ��}~���u#�d����o�>a�ֿ4&��_��0_���^n߶�Af��3Ꞧ˦{ ��Q��GF��n.e��5w۝�đ�}�{�~j)�#��<s
��r���m=I��*��{28�1�v?�mq���"�S�d��m��v2!��zf�m�Ae����Í*���MR8[T��ϝ�T�n���_�-Ԏ� ,>����c��hkt2nٳ{xqA��QƟ�������#Z�J���׾�xlE�-u���3��-�q�HLԔ[�n�vT�p9Q{�Ǟ������i�v�BUe]��!~��E�ㆤ�?q�BP$x���Kw�����넱�q�ѡJ*��ם
�B%����|���ֺl�H��}��X�ioJ}YC�RR-B�q|p(N�#���Aj�(���E:��)�຃����%zq�P`>�t3)�2t#d��%5d&�ݫ�^gD3�͠��0�������L:�6�a:��C1F-��ܑ�.�h�9J�,��J�<�Q�;n�{��p�����T�����v � K�����V�PwU���Ap�b���tT<3	�Tf����&���d%d}��[0��JP�!ܵ�Ƶ�[G���x���x�ĲuE��1=��4��쀋�?���@�^<N���Ũ�/��@�����QE������4��qt��ї*7�ye85ѥ�.�9l��;A��025��b�E�����j.�����2��==�IAj �&���,��wJD_����U��c��mF9��$���X���7�g3�bX{ope�le��.��ښϬ[`���~�Nof�)*�an��A);c�?7;����m�@T��L+v �^W(�O�z�o����v�~ːՍ_��M�O��Y��U8�w��޾�Ѡ\���4�i�����RM@�Y�.j-0��� ��d���V��n�-T�}H�n����gAD$/oӦ.�V�p[=��I����z�dYl���y�89�`R��Z��n]=�c%��P��連��XŶ ��w�M�XO��.���Ԃ���)&4EU������״x	�t�]����}�e2�ZrD�Y�? 95qb�J:T��m�u�7DEe�k�[�9�KY"�D�D�h��#Jl�8�AC �a��q 6��0��Ր��12��Bh�BJ�����zpP�{mJ�Z����v�j�d����jP��{-1t6/�;CKz�k�ЈSI�x� �3�lc��}Y��R|l�IbR1���f$v�|'L�4�:�͐ڙ��!���b>�E~�K��T������i��P�)���"��f<�_셁�p85(�mr�Vj)���� ;�q�#��(9T�n�ۨ�V���[�~�?�Ч�F�~B��!���я�����U���'�Z�EGL���
�`Е͐7`�2��<�A�H	#<E�E'��!gy��oئr����N���IR�0
��-L��J]oJV �L�/��Q+��:Ɇδ��<�n(��d��������|��[n7��d��T�,�Mb@�8��p?)�Ṩ�C(:t }���W��cA�1�9J��+�z��q:�z����aB����qZ�r��\�__՟��]}�'��I&��|bտm��� P���F��x�\;���@�����)�KIk;�X~�,���L	
����ᑬ�f�>Af_#��l5<��VW��1'��Y|���U�Oᬩm3��+*���^FI�a����l%��m��]0�ع��PX��5�
�Ӏ��;5rK꫕����U�-�</�=�k�ƛ�k�&`�$�BlP8�4��G9e�9���k�}֣X�*���gH�:��vЌ�^	��Rq㎘-r+������ҏ9fu��|_Q���t�T�b,j���.Y�ṛvu�)l���A>��7:�PM�'ˌ���	�����ȇ�7�Ќ"���-�82!Wh��ϱ?m��X~]��P���O��+�E� �h�$тK��c'u�*ZVm���P
��^փ�A?���}P����K`�0��v?)�1�D ѾH�RP��+E��b1�J�CZ�m �0���L�#ÐJaW�+sH֯�M�'�OX1s��Ƭ��7QŌk?�E}cl���),����I�f��N����VX^v��%��$`_�Nx���ʐ$��k-���ed�<FX*bVV��e� [QZ�j�k�� �(F�ͥ����|�_u��3Q�̖�,�4a��%9� nb2@�5�G�NoY>ޱ{j��>�:��T���]��Og�n�W�����#PQ�靯6�2��d��+�<�!��A�ɯ޺T������Uw:��L�tTT�򪲪t�*/��+��Y�����"$G��*��0>�.��ӓ%��A4Yr| ��=��e���?�������k�nX��[��H�������xh�"���%{E���5:@���J�\e��� ���%�/�*,���d�E���*!7�����Ao
�Q �HI�>��~�~c��r-���0�̲=V��%�m��V�GETAs��HM0�E����$�s�;�����4 D�1��	>X��!���[������uB'���	ac��"���	�+��%��tj�k2Yy��zo��e.���޵��e��}�����jPP�JB�������%�"��$�~��L�FاȎ��J�_�������-�8��pW����A��d�9�b�+��\!�X�|ԜZ�Mp3J�H��x���匆z1Y�ԃʮ�U�ڶ$���́p'�̈́�}% �c��LK'�6��|ד��d��:�5������e��ΐ���0\�ԥFN��8-z�T�CBJ�Ўh�bI�Bs$3��з�Š���b�qސSJ���s���z^
��J��ƙϱ�Y��ġ��K�F>���a����"�\��KI�G����	�{o�|:��O�댂��<�K�/���}��9Q���	_Ys�Cq�:C��jJ;V��{⬷Akd�8��Un����2K�!a���|mg	Q���)���n�<����4��S�'����5�`�HM��?�>���:��<q���jb_��o=��RE��F�gz�����Vg"}��z��� ��c��6P�b"cl2���P�X�f�,8������0:n�/OM
�����A���cI&G��:����@1�Ow�&����,$��b�TN�i@�_��Ӹ0I���K!�bV=�M���T���͹�(7�AA�a�{I\բ�Hh 5NQ�z�Q���8�A�ia�H�m��.�A�Ǉ��qfRX΢T���K��Ib��Ю:��qyF��#�aSߵEpr���8��)�h� 4���z`d �/�
����֐�?�E����-*�?�M�Ǣ6Ӗ-I��z2.<dh$����=���Bf�1_O`�A)�2Uޫ���롁|�[�s��T��h�k#K��k�!��])^�T�� Xz{�*���H�D�D��o��#�nW�D@��O S�&ruw	����M!�Y��~9Z��6=@ҳ	�R�z>�U`��ba���٭�/�d���
���������u��dv��5��S9��ݪ
"��A����ø_-'��qD��k�_�|�Q�&��z�D �ău���d���#ҽ���X�Sdl+M7O��c�eD���?v�E��=&�:au�G���,����T4�<���4<Xj�(��4��3�
X�[��8u"��7���Œ����v����tqT7&N''� t\�i!H�\�b5�dMi�����9'[��~s{���>)�vdHU�i�e�D��MI��m�LN�Q5����g3�W~��X�y/�5��H?�&$�I����sLll,�KK��?�DL���R\w����7�7:��ˉ:)�x�Uԥh��ؐ��tj�U����u�o-�X�;dk����������۵X�ЁM�kMPE�+t��\I&��Xؓ<;ܽF�����*��@��nT��3䚼�֦'e���8`u�SlX��Ϧ�k�II+t�#Ǽ.oƆ���4Ίr�����x������b�@��q���5�_՜����ۡ�.q��4Xs��W�,9��	�}��$�ecH�b�~�)�B�A����w� ������̵:˹X���IM]�]}rr�KnUqr���@�9�����på�0��w��T�:e]1ǷfCKK��ٝ�� Hߢ�ޓ=�ӀH{P\�E�0d�H	}�k��Dl�4r�K����q*�c}���Sˀ˻dF5���I���
��Bo�iE-��E��D����u����J�v!��zKp���
VB��B�w�g�sp�Tsآ2(k���,�-��>1�{H�Jh2$q'�,�mtP��%������� yS/,�����t<�1���u�T�t��Z�3���*ؽ��Rͧf���a���C�ut�sz!lX�N�҃�	�ʹ�
��3�0^a_%+	,g�5�Q�I���^�@�Ξ�����*���A�&�5��@�5�Һ)��9�H��t�4�fC c�<a���A��D7�+Ċ��0�_kT���L~g����j�̣&-�#O�T��8< ���>�p4��;���$
��;�`��S�l��@�td��s��6z=>��Y�;]o0惞���H ���<��}�  :�o,iC�"���	M��8�B��3�J/������O%�k�d��e?{���������7QX2�ֶ3���uz	�o�7�낋�ϫ�����E�Q�׸q���cZ�-�L�	-ʀ;���A��DP�d����bnD9{�t ��[*��7s��)�Y�_	$��"�5=�Ft�S��,mf��d�̏`[O�U��o=�d�K.�N_�O�o��85��)9�6>2N,׳*��ųL6N�J��uU��gפ�YaVa��7r�^|%N�X�m5�3��Myǚi/�f����p�p���F�q��~����kp�x$p{�M���k)�nG�j�h���L1NYt�&L5�hʫ���ӈR�t�dB{}J	�?�6?���J/��9��$t9k��C�69T�f!u�Q�?q�W��V�����0&�<U����k��r4�$�C'3y�$�]���߻�8t?`kŇ�6�x=l ���{nP#��l�Om��m����u���E�%ŝ�I���O�h>Y!l6�D�"qu6��i9��*��Vi
�:f�(�$�J���:]e�2DCs�[��P���Lď��ϖ:w c@���eF�����n�b�=.��7�ۙ����ͦ�b�c�o��l�iDK���7ޙ|��GŚ��=19�b�p�z�D=��j	�tYg97�p��g'{� &l!�!i��Ń�]��
�{9ڨ$mY�z#���sZ���}=*����0a�Hu�I�cK@�X@D97 M{K�KCJc�f�o�%$!ET��7E�����?v�~gJ�r�1���Ӎ��ΨB��q����sI@$S��k7�*2��$�ϕ�S��c�=d;x��ۂ\�
6�Pg�QN�$�7�ZQd���E����ݴ���FJ�q�X�\��m�I5RPr�Оs)� �������y�	�H�9�5���ñ3�i �S�Z���N\�MM��l�3�� ���T;F@�Z	@M���c�,X�w�g&���p)�V�r�@���P>;ѮC6dH>�|��5_�����~/|�#�rk�y�|�.��g7�RIvһ�^|u���J�Y�͇�dx���C�+�K>���;�S�N�i�-�o*��p��I��W�yA���ЫGD��!0�R�l������S���sv�F�+=+ej�$
�8��1^'��,�@_�tӃ��#.'�/�����j�K`V=�F��m�К�	�z����6��>�WA���>�	�
���Q�>H� ��r,P��BT'T ۤBNa>m�D|�8��~Z�pA�G�j=���Xc����V�;!�Т�����*���C��9N����������K��B��Ye�+�\��ݎ�lW��7��kNO����v�_�d��e=��"	z�cg�jQ:�O�j�ٲ{�o|1�A�
z�@���	�G�f�����d<��>8#�����c7��h��|{������oE���9]�ÿ�������;�w�O ]�𚟌�[	Oڃu����/���V�h%��[E�Z���A�����u����`��U�.q��$���:�C���`�q��a#��^D3�8����Ej~Y�I:�>�3�c�m�V�@��R�褧S�z�,V���hj�0����6���O>nd�{� ����ݙ��.�d44��Y�U9���RGȫ0b�2��PM�Bk�@iq�w�KP����V�s��؎�"/^����Dz $����]�|n^�|ud� ���]Ҋݗ",�=N��B��R�b�e�����m*�#��뷔  �ک� �I���u�H�wg����N-[!ٯ�a��Mѧ�
[	��<V�vEH����5-2ٞ�3ià0�^�$�Gp�'	���d�r�����.A��g��k(�C��_=����4.a�#�4�Q��l#v��"��6��	Դ���j�ɨ�>�d����ĭn ���D���o��2ZyA��[��vw����&{����]�BRw�gU�(����f��gffzsۉJ�v�l�=�VVMhAVt+�ю��h|i'�mGZ�Ipn؂ƕ��hqG)hv�,���}z�W�G�{4�B����C�Q'krE��k=���H�����k V4�o
�\��yZ�κ��t��
՛����CZ�Y��R�kfWk�I�r���#'=zj��u$������(p�$]F���V܅S�4��>�{,9O-=7Z,�'�]���n�爫Q���8��[;�*����o��@�EJ<c��%;��E�b5`�uR:�9S��,H�@ѽ�nj���ߖѹ�U���g���b/��U��2��p/q��2��&�8K���	��4��\���~�H7��^�ݑ��~']�e�V��.���i�',r�����K�te$a��	��&���D�	��Ȱ��Ψ����u�W��R�dw� -������C���
&�ɐ�om��"�J�'��S���+a˗t`ܑgE��6�q����p<*"e���{+_Ua�Y�*�U�*�9M
�$�Ѡ���Y�0�-����@t�8��#WhR��&��������9��a��U.Sx�Q�]��G�I���{%�r����Iq�WJ��"%��6��,��J�g/�6��2��Ws$����H#�$q��%2�����?pJ��fR�PB�:�ƻ��$��ĺ��*8��9wHK���
iw@�d�U5yÄ�}̯�0��3s�N|����;c< ����Y4��˟܋���n�p�
�8P7���^�x����@�>�v��b�b�~�xwrbAP~�˜ިe���"����TF�+ܬ�in;��p?�Ƙ�3T�E����hc���?z��#'()�e�՞νJo
Ȍ���`�(�{M���;�%�5ėL<�+R�O��Ɨz�쌅Z�y\�S�����4^���~�3(����Ѕ�]���p��B�x���	�#��%���B�\K��8�Ɔ�������>�H��k1%KE�pX3ڳ�xH�����L=-�� S��l0���FW�z�>�g�Wʔps`�0V����}�w�L��]�� �`��/ub���d������@'��l�;y򋣏71o
�?Χ`v�C�j�=YN�Q�2�#�ɰ�����=8A�M< ���2��,��P�����6�*��ٚ/ (|B�U���.H����}[Cb�i���UT��$7��X,ۺ��]���.����YH�A=�Ӑ��pU�	�4l��"��׷B`]5w�p�s��2�`��}įY+�[wu�qj��؏�k��@�)q�.+�Th���ܯ>������b�dF��h�IX���p�TW���;�kH?�lš?���s$��q��O	���>�rW~%�,Ӽ��	�$�S�a7���<*�ħI�ʻ����0q��XK6o���2�>>��WR%��v#^,ѩ\��t��,�Ů"��B�k�`�ɗ��)����v�lX:5�$Zր,+\:��V1�g�C4�KgOo ��.���Y��ŧx#7I���pE*­
<$�1��O�M��E��ڹ{?ӿ��Y���!�	�zb	��H��u�ΓW%GG!�'c�rPJ��XT�&Z�E��U�$�B�dNo
}�����j/��8���^p�3�]譾����d8)\�B'��GW�9'x9��d���~rsd�ø�eǀw�;|�vَ�,p��������'%wZЂֹK����p���Qqn=�~��l+έ��N����� ��E���f��ȝH_@eՃB�2)E���쾘"L�[J6�Fb���@s�ulřF����S�_����bBߕ=_r�����~�=�pJwDE��[n6�^�-�Ry+f<q���ܖ
7 ��a�دW�&MH�UOtHK?xP��A�}0�����J�0)\�ꍾkŨc^�HG������ ���VB@���?T��p�c�|�P|tqFك��[_0w���~90�=0��6\��""��[}��؎����;P��T`NZی/6Yr���}�~7z�׵�8����@�bK	�J���M�F����e��BI)��,8�����(m�H6{�Х.`)f��7��Yq9p�1�	Z�'�����yr3c��-�'6a������$��g�P%!j{��m�5B3([��t�\K'x��c���O�jܞX���4�l���"��,�bm���>uJ����e ��,��Z��]�}씢�,��1I<�	��x���p_��ק�hmc�r��;�Q0��vS�~��� ��������OX�[��P޺���teH�w߯sMT�B�W�R�M=�����C���"Nvis�����!�5����/���TƻƊ+��!na���c�X|T4��f��X�*e�U�?��Z������+@��'�ƣ.L�pý�,�����u��R�t�݁/Bi_�]s�c���$��T���_�u2�8��j���|j*�!�{�.����rX�/��DM`Ɉ��������.K�L���cGJ[C������$'�l�Q�� ���,[��i�̗�1ird�(�������d��ˠ�bt�i�_ �P*U�p('��X1�lL����c�}��n64"�g�@Y�fNp�����L?��S�.HL�n<�[�N�#�9QQR���2���y��P��4��8d�V\LE�ݱ�b�E����ÿ����E��W%>Yh:I��7�Ub�Q�����5�6����pR&�Ψ���l ;!MQ�������7��M��`��?���
b�8o�\s� ��XFB4��w�)�����J\����	�?�O8~��@��i��?E�Ȱ���C�	.����QB[鸹
�>pk9~���d���G�H��6��.m���BU5��Z�8��p2�Xl��O�r�7�X�� k��wa7��]���/iO��pZ�99�2�6�f5)�@�π�X!�&	m�ATQS��O�d��edS������B�'(c;^�n;
�/j7���	j=ty��)�D:�F4�⏰F1b+�G����@Q�i�R��on�cٍ6����+�"��Y��i�繟���k�^J���m��B��g<�"�ZO���4��ɨU�ozJ�^���DG��-��r_E�Y Ң̬8�"05��0]Q��1dý�`�[�Nm2k�e��hP��E���ٷo�}��gE����I���[<�����k!�u��%����;^è�9[ڶ�GS��S�"����a�W�06�8q)	�6��.�(¿!+�����
d��N�\$SR�=�Ճ2	�,�T��g<pߜ?v�8��eI/}��=����M��s(�Y�v#E ��1���0PF�����*�fB��@�E�4#s��ߜe-�B�oQ�����v�%{��b���_�,C�� _K���,E5ݶ��E�@q���M6Z*c!��k	�r�]}��	���	$�s�1F��Ϋ"�0+�Μ�f.�|F�ʿ�L��5-�U "�i�"�6��@��|����J׾|}W����$i AjG���qd��=.	����X=
�_D���;V��x�kK��솙�a=+�e�L2�~s�I�m���};L�����P��b�le�c�KbPjq��ܩ���[9&�%��l<�t.BJqX�_*O�T���>�Fa)뇑��\یr3AK�|f����}c�M��L�|B"�aRA���t(�D�@Q`��-E�Ǎ+e���u��P<1����n�N�.#��G}���ә��ML�-��^�H���4U"
�∢5���67����pp���Xꄯ����2n
��O �5�5�6���͒��ʛ��4�tO*�"�=���V�o0*�R}���ꘀ�u����d1�[�9�Yӻ�a�񳕆�3�ab����|3;х$}����>�G�dz���f����TX[�,� 5�ލ��pNK���p�������؎�&�R���0d\�a�q���eK22�S�6��HBuvG>�M�;�����t#)���.�U�C�5f=�7�j�e��Q#g���	��Z��[Ǿ@f_p4���Ģ�fo;w8(�����yk�� �ŶsV�m���}�i�07��L�-e�m,���f�X���Z$-����W�����Zϓ��
� ����<4�k6�+*S��z8a�l��~�8E�"��}@���S�QUR=��s�/��,*D��t�Wϸ�G��ͼ��Z�\U���
�x����E�~7rX�����+k!`���XP�G��͘�'�L���4�e3e�.�@���T�M���^$��:K���rg���d)��&�$�}��`�P�R����7�.�hϙ|���� ��] ˿���D��7Mg/�ď��mՔ��~�a�����t��v<(�q�A�Ї-_eE����e�[�w���fn����'f�֯�l@U4��z�/���b��vt�-/�Xŷ&�E ۶�v������W2M�3��jv��C���E�ߥ�F�1ۜ���u	�m������-�o-����hSH4��a�Xʿ���R
{���h�zU�f|�=D���$üX%���s��}$��SC�JW���k��y���8���[ <.�=Z"���)J�.��Pi�������^����ʩ~��I�T���3L@ϐ!-��:��zE�x�~y���� YCBp9/`=Kg�n|��jM����3�X�x.�'J%���j�3�����Ζ���Yт�	b]�K?�XG 2˟�ֹוF�߈=G�+n�cyq�4Լ�� �6zZ��R��%�jS)2 +��a��$A���Vs����w���em�H��1s�ir�Su=�p>�S�~��E>_�xO�E�HN��N�aܡK�`v~(|�πM6v�&Om�0���m�o&b�a�R�fh�۟f�򜏉`�NF"(
�3�F>	�.�Gr;����{��}�1�}��3�/&�t\�9�
e/�]�h����_�y��m��!C�d
e��6��/��ڈ�-�)��M��&���L��B����K!��e����z|���cZ�)��}R�8ϕ�(7�X�2S �����&�tmo���6���24�,�'#��R�}Q�g�4�[�-����X��r�Q��ٷ�z�8q�8d�;{#[��oc��sz�=��}V]�1�
Q�U)��	�:��O!�q��������v��ںz��v5�m����T�}�SY���#�͇�鐯_Xz>��M6�36cR맡#�"kJ��'6'Z��˃J֟c��ς{��#d6Hk�叡�d�XF��7(K�f�(P,Se��W����){�, ��wgO�G�^l^G޵ro��R%lJ�{r}�VKw� J���}�R���k�v�b{P���(˖aʂ�g�*�o��h�x��X���O����S(�Bz ��gRe��ۦ܀Lm��ltj�g�øoY74l�v�a�jݨ w?���(�_��H���]��J��:�\I� �� �ӊx7��g)���%����%�6��Ĩy�v�26(��J�94g%�7����:$�S��|�:��^��5�	+}�{�Ƹ�G���J�y�ѧ��h������2�P%*x8BF^�P�ˏLA�d��CÛȀ���d2��x��q`Оڋ�{���î,��z�Ä�lj����z���m����y��x�m�F��f�_�'pe��D2�LU@��L;Է !"=�j�7���U�3�w�ݷ���K��#��%c��V^B��b�VH�MI���r72�R��Lبߍ������w��0�$A��ET�;�pU�rh'��v� ��@˧�/�����H�xn���x����b�7�<�ff�uC|Z�m�'~	�1w�������P�Vi���j������(���3:�_�EN�i�IoX2SI#�q�#��8 ǁ3k���n"Ju/�K�U%\I��5�iÜ˖����p��������>&�]���Ǫ��ܵ�H6͠' \���P�`�E���H6)���w(��)&���W%C��Z����^Ñ�.TI؂�쵿�$LDs�U�t�����`�N.W��m��=B�lf�^3���F�1�.r�tCk:��p}V=�J���$k|OkIϻe�T������cF5����<���2@��C��TY��Pr=(x�a�+�c�^�]�S;��y��!|�X�(�`o~��32�H_�
�e#��W��Pѱ����<��4�=̈�o+���D��M�Xsuߪ�ic������s%k��G�V��e����/%U�g��Q̧�k$
�(A�PstҪw'|���H͹`3k�a�)��뗩�2��ޡ-��H2��Ŧ�pq'C�z��cȾ�%d����g���#*-��#d��D���S6�)$�|l��%'+Unڈ_�����t��ɋ��ˠ7����V��;9��{T�5������v
�m��]Jm���<��3��p�7o��}zЄ���������u��#�����r Z1~G��x��?�b�΁ ��nMo+���J���D�a ^i�,�Q�b0��B��Y��g�l ��01.��A��u"<00L�W��aݮu|�W#�5��f�g���j"KhɃ[rP�"��1ū��^x6�?��#�=��IBv�[��8o�7'7	�o�:0N�����2E��\��=���� �*L��&��]a2)s� �F:�.�mT�o�@)��]nˏ������Kj:�o��uD3OZ@����C�?��wL�D+hP7���8
��O�c�LG}��nߪ�x�? �P���{F|���;)���nLq2���va���(X` �9��$VF�W�틨U"2 �G����K��h��Оu�2�y�����#E���%�ᣝ |-��J�8����!K,@���l���^�U�������L��7��e�en�3j!�W��(1������wrD=��ִ
;=�*I�J^m�z��M��|'%���+���'ݕ*��ľ�/���0�6u蹁����uKm@�H�Bex�J�oQA.� �H[<��}��mIa�Vy�{t�W�HG��Ҿ�So�����ߐ��h�TiQX�:�`m�Dp��wWU�ꝗX���9��	e�������=��R�ט�P�1�4��x�IĨ��g�/�*2F~��x�y}B6	;�5�׭��/�F�K<�=�ҁZy���-�9s6�)oˌ�j���`�)�m/M	�f8���4��(�][!t ���W���-���)��Q�b��5�4L58�F���d������0{�&A�=��-���ns萻��
���LO��ˁ�f�/
C��65�Ώ�,p������g*�鶁���3����*�]�T��~��|��%k+� &LG���V�k.����Fn/�}g��5�P�w�	XI14���3��
0_�o�pL)p%���7 {Կh��sײ�#�~2!�Oz &��W��ϼ6�>�VH:W����Ҝ���X�/ _�>���о�-
p���N�`�3�����|���>�5���#�\��=�����~��&!a�n��BC|����k>䃸4�6���@��q�a�\X���7gm���V+�	r|����|~#e/|D�(�R�|A�ad�9Mv���{CU:l5%�<�dz��,�T�Yۚ��$,�ud��g��(uӸ�a�ۑjr�˶�1@0n�g�q���J9��&�zdb�_�g�-t���f�0�`5��!�<<�ͳB�g�Y��Z[�K>�B��h ��"��{�r�}�'���w��J��%�+���T�Xd��%G�m?4�$e1!6#�ן���p��f�+ڨ�P���!�q�;`��Ö_���ѯ.x�ݧ�3�Lst�9_��=���������h��b���x�! D�������>$�� DXn��:���Ư�#A���X���!*
sL� ;O�4�N�[��Tg��!�(�PqVN�p�c�(z�ݠ<�ڼ�]�0�1���,�՚�!��
v�*��y�t��1vp5tO�TusR�ѹ��1G�*"��Z���Y>3�.��}�2�N�$K�kd.�]|�2o<�'ASLδU����Ӽ��:�K0=�(D�Z���'|�1g��4�~����"mO1�,�0��N
��O��eL�+�D'��'?(�d]����A�[�ʘ�o�c���'l��QrAL�ٛ㝪�Ō;�j����R��_�� p��4<�Pcٙ�o�ʚy���!��3��ip�/�XZcm���A��<u�0a�d�ڊ��e��M�N@-ZI�3�U=r��9�DgQ�]���yi���	;~&p_�V$�:���FC���yp��Q ��Y9}�)�G)?�tL?�o�`s�N|y/kz*S�,���E�ұ���W��M:Wr5U�A���H��5����x�޷"��KI��5܎z�}������I������pj^X#�kW#�`�V����A�i�}����ܡ	h�'�(�8��Ʊ�[GEk�j���GJ��̂���ŉ>�5� &x���C���Ƞ��$%LEP
7V�P\Z��
��Ԥ�p���yM��7+��S��Ɵx�ca��MȠ��!z� ��YZ�G�4�'Pa;�#��b�����f�VG�Uנ��# ����&(��x�n��ag�a��y����󁈄�^K:-Z�LU�ohs�z@�D���K|=�`#�����p!���o�[˗Hiżpٮi�i�i]Tm�
���s\^��L;��i�P�2��Ç��o��D�[���zj,`�F�R*;xB2�Z$]�!كF ��)!���4��3&��C, �u�.�K������Y�x5���xI04��VsJ���4RhO��9����0�|��$���YR�ѧG&�)�.��$Շ��b#�V�G̢�%�>�D��E���Et�X��������Y�9ӂ��?3�
�H٢D� TjO	��fްL���|���7��傞OAԋ8~.��5��	�H�/�̪X��vzǨJ���~�lT���&���n;�$Xn��0?A-0����f��2�4)�a�+�n*)x�, m�q��V��V��fT�!Ϭ�7(O���P�F�Q�ϴ/������?��XMw\��ց��!`����i\)�u�������X�.	��oGD���g�(T}��gn�ȕˑ�<��O�����5���`wkԇ��bO2p�ɨ��U���K�>�L���n?F�\ ��mX���SNLǜ��JC����}�������I�D�ψ�O ����`�7�x�Q��yer.3J��Y�U�x<Z�nI �''���[��n,��O��qs�W��W����Cّ��2B���2�(�M)�1`��NGb�	n_:xD�EٹS��7��a��ξ��FRaD���#B����)��15-c,������F�c��'�WX����k���i���B��h���|] �R�����H[Ӷ�Yf�#���fïx�jO��y��1�&0�N�w+ z6�T|��V�P�x�-y}*�APF����i�>/s[>g�9Hf��ޠ��%:2t�ك5M��%<�!#kp�1��2 %��q]�O��.,�)aЃ|�`�2��-{6��]Z�������N��ʁ2י�OŅ?!��<�L�j��@@�TA�q3��*��4�K��M�L}b���֣EO	
<bqC{8	�����v����1�fi}dˌ.	����r�d�=�;X�:U�b�%��_V����G�u�R�K��0��+�m�Ђ9�d��$B��\h��f������5]U3��O���Fxq��o�Ëh�+��%]v�B�6g��x���I�RL���k��o��Sz��-Qb:��t��?� `�$���p8�H1P�.��>׭��/%���)�|5�\�����$�a��g��� s=�*`$�z�, ۪FvA���>Z]�a+���p'Km�iŭ���)�W����I���➐�S(�Xy�Wp�I���� ��~N��
�?�J[r�4�R~�U�cv��s�UP7�g%�R����zh �TR0��LBR!�@��/���aX����M@O�xg�ѮR6�����4�S��SJ �JmBgp$♻��� ;�1�������ӭO�� 9���:*zy2��H��P�T�5��D�L���p6�2#��c���s�m�3�k����1���Iz_Z���Da����J�&���zx��Q�|@/�McX�Ǳޤ]�s!Qzp���� XM�m�ېOH}�A��͝��ݝ$�~Y�I����sF��X
�B^u�@;�:�XD�.�>Q�`8��E�����U&vF��TT��!]�T�IV-�2E�vmg��|��.)�*���5�{c���G1��Õ�S���G���A�i
�A�7�k��TE��/��a���5�"�y@z�?�h2Y.w�d���֍��ʜ�.��%~�]�l���~�z�>6��@Og�2R���oP�PAx���̊�N�w�s�6�߅#J7 ��9�FfԾ�&I�F�Pb�fm�Ӣ��J�n��U���� �q͗_�9{I�T}��߰�T:P�ؙgKԁ�
,q��Sf�4$u���Ҝ���E��;��V2���r�KWt�}�y��J���7R
~�Ism�I���A z��K�+�c߰"����S�M�6��!����o�"���Q)VQo��� :q�JĜz�c�:��v=�( P���p)?�~+x0��]��"ޥ V2�n�x�q{�=�1��Dz���"A����O_�=Qq�m?��̏�`M$7�<���"�y<%�Fb�'[�6�g���.������L`\$��sw#�{���רaHǖBᮣCZ������-��@+cQ����m�8u���t?���:���,t������?=ͺ#�5:I��W^���w��|t�<n�����_Fm��~ka�b9����5��WƟ�`F�jE�^��H���ڬ4R�O��D"��_����4~kj�[5�i�.8~�)��o�0 p��ԫ"�[G4OLi_J�v�s���p'�����6f��mE�m�.[N�N���J�$?y���W9��>�]O���5��XS��I�֘3^;d96��G�U~�6�#��X9rq�}ɤL��v�aayz�K�9�؀1IH8�����4�{�LX�b���?��尲�̟�2���O)í4���Vo�ID_f�J���c�u���;��SVx�gQ�#��?��F���5s��i��i��?�wH�%����u�'���"],�΢Ȏo�A"�l���*apU+�u�,�J&�1�>�n����OO�d��&TM곐r�x�C��.M�{�~͊�1�ҷ��4���{+a���p�͍z��K��x��="��8�
��Vi�fk�<�3��C��ER�/�Y��N�[�6�]w\_-j�|�pr��j��]�!]Y�Q�l_�Z�����K�i��u��P(�\�E�|��G>D㰾F���s���a��?�dҲ^�
��,OgU�M=pP�yi��[W���'�'���lY����3^�H9�zї^��� &!����
Zq����L�iY��| go�7FlI*G1(�O@�?�La0$����ֈ+v���i=�ou��4�m%4'z}%�2)(���|I��~t�&���2��m��D@�N�E��Nu�TUV�Z�|���O�Ge�G���η��	��3h4Q@8�_��遼m���}��e�}�gB����=�{��f����n1���~�f���?�$C�� �8j�M�%���4,!��ʺx�c�|�ؑ��*��_�ʔ~wf�4�.�h !�����~���Y��� ?�٫��Z���d�D������(d�YlB��ʵcI�Ҳ�K����jk-d[��^�$ �@X�Y<���2��\��H����1���pۄE��SY!uE�{~�n�DL!�AK�1!�)�Xx��Q�,nB�X�M����Pa[Ml,��'��9{�<t�'�s/	�xj�"����}v��!,SH���@jXBz��=�K��1b09�H�n
U ��G�6'$\�����iw8[�N�T�h٬'�"�q�t�ܞ��p7����М-A�Xlh�/8�gz�&�%R�<��d�Q���i?Jj/� ��Mb�< G|.����{EoS�8��3>�;wBaQ�V���|6_�6��BMp1�J�T;Gz ��#�� ������0L��J��+�PZ�B��G(FؓY|$$�(�t7���m�<Ap�j��vI�9���5a�;�?Fq��ѻHL�uZ�Kw�y��l_v��Ţwnn&m�ʓ�-b�2#�T1wD����HirL�U�z�Xu�W�� �³m��2t�t�Y]��|����(&�iT_�1�?�#:
V�Rft�;���1c!¶g�R���&��y{��ו��+m��n`��A�(���N�I�#6��B/��_�b��W�-���$�t���h�
�n�ݏy��wJ}��7���o�i��P-gƀ��-�x�7��d6k�w��{/�6����R�3j��i��1By�-���+J}�"�����Q�֧����N�_~�3�=���b�o����T���r*�*Ѩ�*t�X��M�����r�Kts�:f�}�_i�~IeW�o�nútL�\���k��e�3�h����~����4� ��@>K�C��bPI�a��x�B\N�_�-��[�oi�]ÊX�I�x��\���j;��s���-Okl�+���UkMoxeCO�Ɔ�[���%���t^Y�5N%P�G"r��Ek!��i��a����ɈD�Ua������٥m�m��lL�b�qi1�
`�ld^y=�v?)l�7x�Z�W��!I@Ŝ���l2����ǻ��c�" ��9r��*]=l������\^'\���dW��������y�u���Ѩa��"�e4��)������n�_��"5&�دբ`�HL��hR}ǩ:����+qp2X�R�y��8	mvW���L�ژNG`9e0��.��.I���:g! ����QJ]�su�CN{�nG�*[(��]ا��������x�� \r�(��6/�= 6:���IQ-��u�O͞E����B��Ed�d�MV3�#]��N���.�H����+_S���A�i䆒�ս����W�l\��&Ɂf�K?������T,)�4DCu$CnR�)��um��A���YRpg��" ��+��ܐR�BR����GIq)\)Lnp�<�v�#]�VG.�U�!kc x|��^r��/Iz����&��S��ʢ��E�,�x�r��R}�4���2uY(�}�Gb��R8K��۝�Ӥ]L-�z�Y!�<���W�iy��q՘����Qw���#YQ7u�Z� D��
���A�d��V�Ƃ*��f�I��Ț��k����j"��pv��Gܔ2�"���\�v��S�>=���!�ST��_߆�>=m8��!��j�r�YR�8<<9J�PZ�x�S����˭vЖQ\)
F�(��>8Ӄ5�J��~t߿�r d�u}&��4��/��a�@ Sh3�9	 $U���F?}���Y�����
z��TZ��E/���v��O��)�-���7#$m��I������հ�y*�o��0з^BQlz�#�N�!MuņO�.�A��ƳK ���]��Ss��ˆ h���S��R�c���>�+�Ԙ�b1�{��T:|��ɣ��M3g�󐰐uZ�
]���N.������%.
���P�ג�C�ћ����vX��E��T�u}�2�˰����b@�C�Z&0�w �*e(�dRmO�!,�3N,��;r����sqY�@�~�L���.!th	�iS��vW��+-��#�r�d��|bݒB��[���%��K&
1� /�ا�E�<�`E�
"3�i�D���^o?�DvF<S�������_�Q-*T)��u�!�譲a�Q�����)!Xn���� �ˁ�#�JG� ^�)����Q� ���{<��gT��2�6:��i�M�I!o\��< rDpoQ���?�nI���>�D,_�a=��-��U�`s�����KI��!f��ǭ>�&�6|�X_7 ��B��u"S&�z,�7��3�y>�c{?��ݨ�Xf��Bb�ţ���[�%�������B�?���V�m<�4ۊ��u��_r�����j��,	K�:t�3�u�Nd�[��Zv�{���E��4����1��/����3��'�YZ��$ad'�v�߆	$<�=��`���;%Q���``�U~e1���t���d�1��
0%�r�e��MDu���g��������}3��@�}˵mN�$�aR��?��Ԅwj>(?h>h�b|��t�-0#s�Q��n{��w��6�0�<�܁�P#�Y	ՁK���8�Q��t�9��/x����Q?f��T���d\'H7��a���g�hd�}�<?�q��K�l����X��	�k�I�:�_��� 3ӟ��G�dQ�0o�S��H�5�f�ݬY{�u�	L�((�3?��6��ס�6����3���=����׿�tq�(����Ԕbq��8�WGm"��	�������u�).��ߥAj$�k<e�艴n]�g4�H��D�H/�q�.��lIt��!"��+g7/���V;���Puyvة��M�qX�J�}�Zlr.4�D�	�t���aι?E�&a�h�6p��M�(�ج��\	$�͐��F�'��X6���k�ּ�P��3�wW�� �Re��$�l���[��6��|�q���%�7휻�|��!�����8�иt����~B��L�ϳr
�.�7/�Q���W���� �;�q�����w���}:���%)�oM�gt4�LO��=��ƅ���;;�j�k[���s)r�.K��p��I������C)�0Tu#嵝�����t��ۆ�U�"�o�F�a8�_�T`����K2#�7Ȧ�)�Ƙ!�r#OP9J�Q$�6��JQ|�S�kA�5��n"��[mp����X}eW~8�����V�uw��|� �ɐ��5s^7{�<�ѵ��lA��N��K[[N<�$Տ����5���� '���t��, ��
S#���!�T�Ao�a�s��DH���դ<�?��C{�G�_��Qӆ'�I9 w&I��
��&&˿ޫ��2I(��@�:q�8e�ڌ��5�����XAzM�iBG�Xe��"���O=�2�{�(m�I�k^}),*	D�flw�C&�J��l-4]�J��˰Y�ʳÏ@���@%�c�-O(a��U�_`mm�4�(ّܯ6SC����얫�}c�e�bWuq:�Q[����	RD~���|I|%^|��J�}H��k�G�W\�`�ۂ�'	���A��-i$c(�"���+e��e�[o�9nr�ү�����W	�t�Dn�}qSqw}���>�N�)W7b����\�)}��&�Fh��HQ]~�:yaV����ߢ�[H|⊞>༫�O�u������F�>���~Z��v��A�j�:�5�R.�(��:T�r���}�Ϲ�Nl��
A�~�u*��d�/���l��ݪu�ЇA,H��y՞�\@ާ����5f�э:�y�f�D��_��-M�5�ݑĔ����V����!��~��)��&�N�����v���������H4�H��r��:r�[iM�Ȩ�W����
����Mx��M@N�MgC���7�׶���_)������<����������5�/��؏ #%E�"9� glMֈ����PU~��advү"�rw1.��]�X3�:��0�uվ�p���fQH̖�;2�Q|��p���A�1O||C���.��iۭS�5uV������9	{�4�Fr��o�}���YԎ��>hf���j_"��)��S�z�|vq�����Pn�6^6��qv)��yk�ĝn|:j�7}C������d�Tf���7���"V�0��*x�m����6�'
Tr��J[��еp��C(���`����!c'�%�&�M�Ȥ�KZ�2',[�*]�����v\�g~zH$�3=5���\�{�Y&�X�ڰ���@MK�x��>�NTw�pҠb�����ݜ��Z8��
������)�G��G��Ɵh��2�
���8��}<X��ͳ�Y�,�&韁�ϐ�ѢhQ�R�8�:�		���4�QI]U���ĪV+�\Ywr��B��}Ξ����${��(>kh�e2���JbQğ.g?EܿS\g���b?�*�_ɫ�7�!���f�!rh�i>��;(tvL����c��ĵ�~t��ݣ�¨a�*#͸�~ih��5�7�MjQh�WPjq�r0�!�p	r��gW���$5�6����@&tM����f�����^������?i+~�
��d������g��3�rf�r\�V�|\���>ґ���|��F�+��Vx��6���3��bàE���Զ���3�:���9I;@� �J�������s��bĶ�mq]L���$�t���4��%!�xA�do8�����@�ů!P�a\M�.qՠ�"^f�j��":������m�$}I�AN|艧�P۱XJɭ�����
��p�K�@�1:7`t=�f֐S�w��7�zuR�����)~� �s�t�����#��F�CqiI��v����s�TIGqS�e|dTk��K<����u�n��T�탁�^Y����ԙ���h�Z�j�a��w	��#�tu���ʨ�=��a��`F(tQ,�fV�S�
n� � ��/^�^?�+�c�L��[�f��5��N���bMBC�a�o�?=O��!5����_�
�6�d���Νr?��;��%��4��f/�p�ޅ�A[��H;�{7�;�S�\��z��m�ݸ�?�1�E��^7��e���!p;|o
�t��8ӚHE�f�U���3y����G�U�P傶�܆��/~H�b5��$��;�-��$\�!x��b��� rPϟ������Ux�i���A8�T���9��=�Th���ÃJy��/�{�	�����@ɉ�P���+��hWZ�����0&��]�X42��i�f�D��Ӣ���XG���ؖ�S��.���"L�p��HS֝��}�ʫE������L���E5�UEAja!%J���s`E7Yj�Vn��U
@!��� ���}���vT:VRGD�����+3tX�FUzji��d7ͻ���w3��ydȰ�e��pB�U)�$��V�wC|�@T����Š֝:���j�㿶�=/+�:�������qg���g��uN�>V�뒳��%�F�|Nq嗅X�� �p��m�+�سE>�+��6[e�pr�z�HB[�V��S�o��Oͬ��?KeQְ��,�x�N�(���?k��/L~���	
:^<�t
��J
�[+@�N��3�jz��b˖�6 0V���ʼ���/-��G�.�\�&��!Z�������n*g�g�J[V�?�m�hZ�(�[(�w��SOc2�~�Q��ڛiPl�e�#�����).P��D�)l�K�4"���C�k�^JG0_X�P&T�Ku��@��IN�K�P H���+�a}�h	�m���a�#�xEt���.�'� ��ls��z|0�.�=+��Iy���Ï��&/�0EH�����,4
������Uf1K�`I�<�@5��]?����� cM���o(�R΂�(���� }��da����1������B��������A֒d�%�F.�v��$p�bө�H�J��;	"� ��9�B��qq��I)�|���}{��A��I<��&���c#g$]A�8�w8Qw�uad=����	�>���挆/��Ĳ����|���� �X�z�;Kv��Y5����0�i���5x��;8s�I!�|m(-ጯ�֍<���B_OM�c��J-`���q�����7�[���jQoc!kx��$@�u���0R�:�̥h-�Ic;���z�GF�u����»���Tz"��ٰ��А���/��9@�Ԯ���?ֿ?��jVo��_p���$�|Z�L%V+����j��-�I۱$���9�7�i<�� �Yv'�qզ=?	ԇ�(�F�aF:(�{�%�fF��A��_\]�ʯ�(����1�`�A���ăUy�G�9!�����:v�hUM/#��9��c[�5�\�5��RJ����"E��Ӳb�r�B�=�~N��y�	<��J��е��U���b�e�� ū���^̊�$ ��ll����֬g��iF5נ.Z�ј̑ �[�#�����(��<��^�<�e�L���v���w'��F�4�9I�̇�?M?�ޮw�pQ��`ބzO��=ܪ�oCc���ɻ1T( ɟ=�h��A�C�d��P������x:d�����v�6H.�o�\�|��Q]�3=jE�w���i��ddy���/rǁff�=M����f�~LL�:4��G��|��dUN�x�i.�^j�]Q�q���"���Ԧ�%s��tF�qP|����4b2e�����E�z����6k���
T�Z�IR��Ȅ��v�f$�+�.����ŉl���X�&��ur��7Xڕ���2��73��T�۝B����U���q�z�W~@�d��6 lt�b�ã��� �dw��S��x�_r��(����w$�:�>א����w�v*��/Y�1,�f��/�KcG�b3����k��Y ��(�"P�P;Aל��m���B�Q)�
�]%�Y�E�y&�D��4ԍ�R�% �� ��Ia����Bs\�&(�S�ٱ
�t���x�a'g���������κl\ߕ�t���\xMJ}A"h<���.�k�u����Z�3�)0	#�7<�8E�*x�Y�kȡ�$II7�����Č^G;RB�
�롴z�P�T�2iͦ�w�qVkߥS:M�}W�jͤ�e-.!Њ͘����>2��1�� �P��42^�]�]��dp��v���ձ���\��#wE����"};��@~E��i�S)���o[\|�n:ےj�0ج�ӓ���Z<'�#��4c��J�1_��ldG����i����ot/vhs�p�7��V��*B�i01��]�Ӯ���k�x�Sf���A�m�CY7Xww�޳��P��������
3��ɮ�U�����h�4���'m��t��:����;���Y͙���� WGk��)��dL6^^ ������_O�ר�o�_�L�҉Z��RV�%�R��U^ʛe�:_!8=u�~�Q[�qˤmle�o�3j����KK�r7nGo��}Cڹ�-���+�S���C�Fm}�V� П�2�#����p��D$ܳ�k��O7W�H�*���m���S�^����IZ������`���CT�!���Z�=���K��#@��[.}�)�w��;o�lOF�	��8k4�%s���j��H�<y�DK����d�|~�ںh�y�W	��'fj {���7G�+�@_�z	#�̒�q��6�ѧ�̪��ŦB�Og^B5�j�'"�؝:k�'��3���di���dT`��E�\�#	�ԙÊbH�Hk�]Yם��(����N�ԣ��W�� D�q�PFs�i]�[P�.1�"�s�i�ے/~�vo<v>s�w�ܾw�>75���D? >)eٔ�W�%��<w���YL�װ,�(5Q�o�׆�� :��J!]"^�n�fdH�sLq�fcU���^ޕ���VL&�,�/�0��W�����n��T����"�9�d�*���7���fE��bw��<�3�~!���`�@��N�2�~�3ñp�a�ֺ�úߩ������<���7$�N�7���R�7�?Xd��4y
�5��z�,��P��h	>0�67u0ˈ�I�rhלA����s`���8)֔���$k��m)�wOmLI��U�_E	�nya��
��u:�ZY�z���f���֣L�1�4{&�]�tI#���h�|I�q���0�w���tV�C9�7//�	�'����΄��c���9-�?�o�p���"��Ԑ���e���]�Q3�eGme�+1��������'���-�M������Z�ESD��a��l�N��-��uB��LZ��	֫Fo� 
�A��N��������`u��A]])3poS`r��5I���>��"��p1��x�@ǰ����с�"ʣ��5�#cd,��-���+�� �6��a(G�F�:^��7Sg�K�|�z�m�]�T����p��cX+]M�"N��#&y�cL��9�e��R�1Wx۔�� ��&�C�o}��	>eh3z�K��g��[�jc��u�*j2�����^�w�o%ĚC��L%�|v:�>H�l�ɪF�#I�}(#b�|t��3yH	����+r�$&���f�b"W�R�(�6�!�X���s�N��-"2��+)P�����`$�M�z�A�rj�u����]�!g��d�Y�-t�؃H�Y��z��6�iݕ�)p�Vb�R1i)ۈ7�=�mv�m��'[;���g���켡�DF+��V��^Θ��̚�ݝa��ە܀��+G��������(����9{�A:��%�����1�غW�,�c��kt�H�)d<@���p����B��#"��tOeyf�M	��%O�$�x������"����bwD���y!7�ڍ�C0:��H8�T���S㺃�(ʫ{�������,���PS�� �k��r�&�*l�Ʃ��A��ߛ&�3$('��<�7<8�`�<���\�w�l��4���&<�I��dS���z�NYL�nt7r��h���4���4�G�Ks��C��VJ��	5
�YO}��f�P|������h�]i����Z"��$h�$@�<���+D�V��j������q��w�U�ƀ�cyI�$�'%�1�<"��X{�O,�@ג�� ݳ�=O�1����u�mx������S�z��-(e���jqfѣU=�yوjY ���P�ɤ����م�R�G��- �@V�D��cjT�9ͩ� ��1��������>����Y��OÑ�!�o1��,̽�Lf�R��i�w|��?�w_�u��ڡ*�{���+�q����	U�ZZ@q�gN��A'KGS���*����+[ͮE}��pG�^t��=la���FHf.���j�s_ڔC�7S���%���bc���h�A�lT����A	K�t9����´�Z �w^e�)��2�Q	�a��Q;;����E��\;S Uޖ=i�@�ɉ����=?e���?�U����ф9���&GM7���~���mE��Bc�.i�!<��"z�O�i뢊��m�:��gQ\����sԍ�Ԧos�@��٬�ځjiGv���KY������f�^�1�D�y^Rw'�.�C��;k?��F�	zH�@?�@f�d@����F��2��H����	��~ш���Z����e�\�2&�m�K@1J�
"e�z�������&\��W;�]���g�'z�e���D�u��PK��,RL��^p�=�����ra�\��*��z��q�f&(*��l�Ɔ�$�W[�.�X_�З44j��
��$a Aܿ��$"��z3"��@ߪQ?Q�����P�c��ɻ�7r��t�1rʽPl]�n��qԡ�1 ��|S*k;o�E�^���ʢ�N֢��]�@��O��Ƌ |�Q%�K�(�.�6	�@ \�r
5�z"����s}g	E�@��F��X�2�/�]�7��+����nV��Aj���C���	{��e|�?�D��ǼF1ɼ�8�uW�V����X�:���Oc�w{��V��� o����'*;�h��GG  �f{�K[�Q7�#
okN�˺b�Tu�P(A�P)Ʀ�n-�}fe���`��+{��jsə@~^�(�
\B|�>޳�{��uMH��bESqgU�!��L�fK��8�G��dfcEC��С���m�Wy\w�S��O،~�=I���!߽���sU_8�{a:�b�a)�leH�R�G�`�;?Kƥ���๺��*@%%�(�\R�.v�R�t
�� �8SH������8o������-5��(�U���i=�jq8!L���h����<�����Si�ٌ��9�|o���<����ˊ�r9߇ꃣ���\%֎Ԙ�Q���rH�_M���G�z��E�l���^r���B&G��M�����"*��7�*���ĉ��Jҏ���/0�<�y��x�6� �h�^�����U�mo�K�ԷJ��C=2�Q����`h��r��������t.��2TiZ�a�^2���t����S���/�I��Ƅ�0稛�	�8���i�@��]哐d Cw��2<D&�yI0�Ļs0�)����Q5�s~��eSG���V�����?4�qr,N{T�P�_6��Ḧ���*���8up�6 %)k��i�Uys(�Xk��M�^���6e�^[��<�ư~F�`���a�޶�-I������5v��	\���"W�� ż%�c�츥L�&��p��$:���6Ŋ4�?6_��)�!��}�PA��o+Y��E�~���n�Q��=n,I���h�C��Un�//x�*�O�s*¹� �;�Y&+5yO:�8�k���9(��Cʗ�t��c��f�:�}�/���zMv�?yGR��
��F9^�e���m/������5�Gvu_�X���
�Ƀ�'Y�=��:��C�q��'��e�o�4>[I��I��O��j���-=4��S��N���2!%�z��F�����Ыs��ͫ���/��?���_+���b�t��8_D���V��ȃ���U��4=? N�]j#�c�y=�n�T���Ά���=[ b�_��m�7�e����*Q<Y�\S��7�Ɇ���rs�=�1�S�oD"��3pk��6BEW�~��=D�3�����M������R8��2f>�p�v�>"��<Ř�Dl�- w7�̳JYqn���[��"�nΒ�=�y�8��r��(l�[x����Q�*ddYse��Ӆ߉��<�a�QM2�YA�V,�Kk��	/"��C}� ����R���F�'Is�o��$~��K��$.v�6����[/4e)0�c!}�ڑ,��͜fa9L
`���w��p1?)d�"!�t@�k�V{��]�4�Lh��i~%���IzC�p�e5�V�DXg4I��_±��F`^����>l����q�^��ir��'`�	���5�8���y��8_=uZӈ䁼g�~do!��J�|�pQ9��C��Փ�[MBGA��ܽ^~��Nic�n��?&BԖW]7��G�ǻsc�n���X
�.�>�&���\Ï��be\�@	pЍ(�e6ޡ¹z�}"~�-n�3k��?1v���5�}�Be��A�ĿlF>�z�����L�(Nt��S�o�)`+
���D�C��,��s;�u���.�!�k����BZ��s_�N�;��U$a"��TS���L����҃v�Di�ڃ�z���zG�M��c�~��Ǳ&lN��E������e��}'�V�V:!)rxp6�$ D/].��u�K8��0���?�<D�=4h�tȃ�������K��"R�޾$�Lؘ�n�a�2� �����А?����c�Ρ����(��-@/%��_�q__�r��u4��
C�ue?2G��_�%V���e�^tK�j4<,�ԟ�w�q�_S`{��]�Q�`��ח'@~]<J��w��ʫ�%(:��ҫ��k
ϋ����콩,��k�rz�n��V�x�^�	�q�m����ub���S���t��@���6�%E�9�1Py�l����_�ƙCx��D\���t��p�C�*�U�у��ҋ�v�-���!�j��j'�梮P���_���H�(]�!Z�ə���[g�:��p����腫DAڋ�lॉAd����>���;>�o��F#[�T]8`r_�$A���jt(Æ�o�S����p�:M�\)�#�Ѥ����O�i"�j���cRswe�
Y�ԖtД�����Ĺ�k�P/�`h��+PUW�� �r�9 fh{�Í��������Xc�)�Nm?��w�_���d�Šp�wv��|���D_�g2���:[��^&D�=ޕ𰃍�k2�tį��(=ξ�q����(��d;�zcC�1�撋��qphH]O��X<��`>� ��Lf_V<���!Hz�p����׎�s��#�����1N�[l����Nxg�Z���Y��)-i�z��nA��ϟ,O�¥a����{������
9Z�S}�������[�m?���/���Պ㤑�����$lf�f��l�D���Pz���ra�v�)�z�MC�]�&H>��P<�m��Oh��I���طd��3E�T����'_p�����L�ӑ�W	��6� �ͱO9����tzow���*"���%TW�䀓�n���"W���N�I�@T5{O~�(Q8gV�d,��q��������Qmn_��.�3��x�k�_�!"�>d������֥>ʣu���OVs�3zM�2����4��'���QP���Bw�~�����+\]d��u��䅞Ԋ}Q�g3�&㐢��1]�8P�IS)F��'3�4*������Tˊ������;��^����|?oO4�S{<�&p���N��[��r�o!�el�� ؗ8����BkN}uz��0$:c| `W�O�ोL�2}Rcށ�v�7�68��/!;T�I+�&�[뿋��I����H��~RX�)FDJ�6Fw�K�+�lJ���$8j�v���/O��9c�����v%��8�o�_�|~�2cUI�ufF������������@:�Y���z:�mZ[I.ǩҏ�#�O'~}��b�2[�n�n��ŭ�<�x#*���X��XxT��#��~im�%��X��'i���9�Ə�"�l��pDL��U[=�%$�D�i9�k۫ݚu��BA&��T	�n;F���;��#�4��R4�L�!B���,G�/���u}F0)~�����yI4 �+��.�H�xtRg��M2T@�Ү���b����,�,Df����(��`�f�s�z?����aK�20��P�L��>��K�O��6P�g�#f!�V��7����+�cN/�B��������wT�.a�ʢ�$��P!k�H�M��8}�d�=o��{�*]oC�7Uz����N�ץru��ٜ��ܑ�-x.�����w���`�������G��O�&Ն��M?�u�T���J��]-)׉Q�wDY�	? /�+j�Uó]���I���.��,>|�,��0�����o�R2\eۘ�_���*����;.yL,����Eyv‑��M<�nTZ�4`�kCp�l@�73�v�U��7h	�f����p�&p�Y#z*��T���ݳ��e56wL��7z�_v2A�Gr���q���Yu��~��t�{RVk�*!�*�DF�c!p��.g��Q����=[u� �!7�ܾ���+9N�V �/0*�j�pܥ�1r��e�I'���{#=Ж�ґK 8����o�T�V�}��^%�H2�h=.�[-j�w���F�>�8�w���{2U�n�C�F��84����04	3pƋ}E�����\f�O���܇;B�c)rq?��&W� �W���a�>��@t��~�h�W�_* �!P��B�G�vuI���j.�]�ԍ�S_`$��X�%aPe�mD�.h8!(�
���)W�t��/��n���=��T��O��.2�A#����3��8η�len��Q�ŕ~�
O�g�`�p�Ҡ1���A��Q���G��>��c��X���l�=x^�S6�u��:Qc�v��$����\]b���a9��� �%yۈʫ�A�`���q�q���:}Cǹ�l�|i�?=HM��h�,�n�S%|���n�R<*�o�;o�*��:a�3 ]��2[���?�:� �s�襞���k)�e��^U�1�I
�!!k�`��Uv7��@�N����w��&���J`�%0߼�_���!��?���z���?%�>���t��3�<fQ�~�v`ϗ��Lwx�z�\+�{N��a�C�:�-E���Hwy1��Y���1u���^=EBt1D,��T<1ʑ���,]�Y*�����l#��0Z��<���lv��gy�G����m�X7����^Kc]&�W�ȗG��uLnzb���6�=�:H��T�F��'�5���9��l�����������8��~�S#���Qݧ_Hs�_Sfc&��s �zN�>��5ݑ`=-��ጮs���m5��lEq��6@��_���|5� Ax}�"n�1�lBQ��Ͷ=���'0���{ق�DƋ�'>��rA܌��Qg~�*iW�\�F�r�~G�ڿ8����)�;�6p��P���x�v.O��Qӧ�W�ܜ���+��2q�"�S�=.{:��UV�'<���t/!b��!׀��e��#�.�oJ�dO�oyk�����j��C�3f��F+(�9��؎���LE*�o]��n�s��a�_���W���o�yw'��2�]P�����q�.1Em���*; ��;��W�\[�ca�,���&d�8��Mޙ�t���HJ��7�i�Vc텃���II�W��U�LW�"tR8CN�8�������$�E�s~^����>� ����=��Q_!�<[ƔȈ"��FQИYL$5˞ƞ�I8�|�U���8laݩ��5��@pG�&���$l$R�gݺ(c���A�h����鞔�|$����K~G���j��F�.)�0u�Q�z��# �RI�U���%���	�w�h����������
$�;�Y�������G��(٥�8�k:2�s0@:�C��g±gE���p̑YG1r�����rh
����������C-��F�}�a�N����w���}и#d@��O2�Z�oQY�z���v���}#��K�(�ܵ��ًYf��Vp���*ژ����������k{(�_�A��@���}�W��7)��U�9�s���˝�1f������'�ͣtw>�z֊y6P�м��c^мj�*r㛧�<��s�\z�8-r�<��
.`*�i<1����q�ri2� �uSB[��1�Y�
�dtx0/j��.7F�~�	��qT���3�6L�������
�HKYC�Vd�:j��F�ajٓs5)��j=_�Iu��"��-����7	�w��thɻ#Vo4:�$�@�r5z�Sں�V�Iz�a�*�Fj4�%�P4��,��rfh����Nf�6⳩��� �ܳ��l��|IT\{��\����L������S*QʑJo��G��/R>���$��}4�^f��v<�I�8���8o����E?5���[w�<��P��Ĝ7&������ ��_����8�#���1��5�⻹@1��PBgf@g�H:X���� G]ˉ�ѭ����5�F|n�N'tqp�rH����!�����
۴��l���G�e�&�7�6 �~�1�R|���:�����)�9�~%ΐ�z��|rO�bGR��p|��2P���,���jg�WP8	H�Q�o�U�~j(�I��N
���A��z���؄�t�j6�V���	y�u�'�n���C�G�pww������j��/H�q�)���5Oa�Z��l�FK�(�і�'�6�6��b
�u��F�����t��O��6���;Ctax�tj�"���p�i�nyb�
�9U�n����Mp\r���%'fS�n����f�0�T�HG��ޮ۱��C��� �â�<�i��pq�1�2\xf�Sz,@2�"�3��AM�C}�z7��Q�tN����ꦫ�$��2��M}~ε;��3{�����	�U�h��D��+j��;�y/{$ ���1�X�=��(�{GF�=dG��	��XM0������2�\�ad�
P{�G략o���N~G��vP�!}��D�7sm�ߒ&ת�/`�#�]�!�&QbC��|�ڊh�9�{j�	�#`��Mcx��������� D.���;��$�cy��;2�b82���v&7��~u$�Jd�K��P�)@F�.�H�!|zH���rm2,W��C�g�k�ug���4���&�7;,�� ��9��:4�i���z�Ob��7�^�Y,���(�Y���Jjx�9�l�V�#�����U.$��a�^^@�]�9Z��Zu���@��g#�G��Y��gxKg	���,1>� "f��_բ���B ��̳B�_ќ�#��AXr�w���0�;��$坲}�7�ex ��X�v=��/LU4���V^�U�|ӝ(�OD�0����H��M�C���K|L#+�ÍN��wù����Pa��?pF�9M�ڢ�t�Q�}� ��4ll6o6��S[!�F�۞��4Yk���t%o�����Gaa�,��t	��|O��3���������mh�����9�*��9RT�L�n�*������-~�DId���C�J��2u�w�M�,Z����F�ŗ6q����q�|�{LA�h^pX-	����+E��,r5�X����	fO%>�[�h���
̍:���/G�NX�����%�eK�=%'+T��1��J��'3�!Y�%
�!��3U����vܞ�-�:{���D_m̾>B2�
�u�Niv�M*H���h��/�/��,��]u�����_����4��<� M=#�ݪ2ъ���=� "���.���$�~����gM�07 �����s�`��Mծ �?#��а\�H������ۼ$�H�Y�+�y�G���@�D�aN �x���w��An�gSiW���Xn��`C䎉$�������#r�H.-�YՁ$2`ҕ("���)P���ʙ6��[�Dim����@�H�G_Y
��#7�*�YN�+��R����w��P��1h�/x�n?��:�4si��� ����o�B���{;z}�Ѝ6ب� 2D���NW<�3J�jq�/)6ӱ8]z�^���Ӕt�qs�x��Jx��lp@�u0(d�g�?��Bh���2F�Y7[��s�|B��I�ށ�᠗1�:��ih��@��R��A�J�>�>A���"q���>v��47�ã&�O]�j�O��"�2l�v��{J��K�'j�A.��փ���' c,���wTQ��#1�m*�0G����I&~_�wp+����S�V�x�x������	��uf4�i^U?Q�g��,GN��΀��#��'�|y���=e��z�k��kq���X�X��Я	��c��;-B���WmkY��W�UB�w�SՕm�F>ve��>YU�JV8O��B�
��@?0���`��F���f	7�l�����9���{��\'�]0Z@P�U�"�I���)4d-|c}\���{��#��=���׼��Ŵ?��Q�	�~~!���j�b�2�p/��>v�Y#`)��1\�nJ(�Xe����j&�P 7����{��~H��B����;��ePH�'~�eIQ86�,Nh��|"-�s��e����zYl�s���\�����e*�oY2h������c�f���<�M��V��j��H��c� �f�e_݃)�D�q�;��|@d����c���@Թ
k������;`�T��Uʉ���w�;v!�D�C��i��ٱ=��s�RQ��KA$7�'��9II���>�[	<29rS�˨�!��j��?t��Dj��N��~Q?f�x�NM}��!����d4��y
"A(��=@�؅y'Y1�~՞�;�زK�ޥ1�C�*��%'ǣ �g����6wp6�Uصy�f?Df��l��Vp�O/�Y���d�����9�Lz���q��_�Q���|Za�l)64K��&$ #Mu�mN�kK����Q�j)U�Jd�藢#�|)ٚ�a��Uc��km�jݐW^`�j�J3噫��.H�����w��19'6�r��ZK`���虷(��d�\"�NF�v��z�gy�̭j��2��25��\��1����3/��s0H��a��K^�GG&y]$�C��ƃ{�]U�S&̎@v�Ֆ�e�B?����wxT	q�s��M��yاU����2B4ߌ��r�{))�D|}�������w-��3�J�e�wВ:�U�	� ���Z�����i�J^'r����E�niyIo��]�7�����iWڈL�c����1��*�c���h�:�kj;E[z��<��!P�uFb(`PC��B* �vl+���Y&���
тx�˷o�zf{j%|[&��L6�rT"Fe/�YNI��A:�a
�l�JC*��-����)���D��QԊ$`��a5���nӧB; ��R��U�#��ˇ�`�dq{F$� Z��`�לK��u#�>��c
;@@�)��kS\�;������`��z�K$�I��Z��B�%�aX�NZ'0x٥uqQziu�ćp<��~��-�!{$Ex���.�Y���a�'�MB��b��Ɏ1Dבҁ)�j�`�;�F]�Y���vxh�޾t����Z����&��>�V����M�%�m��0 �L��镴U��O�����4�y��~���#a	A���@D���jE��u'	=��#��	�+sxLu��-Fs���wI��#��g��ԏ�	r����ܣ·7�e�	�R>�(E)$q����0�<����N q���}GC_�ν���j�e��`����f��xW�7��0�b�ad�һ:,�f��s�խ�[iݾORT�Ț�tgroc�~�մNȰ���
�h�2Y(��5q1����?Fm�-0���9~kL>��`�V��6���B��YP�[���R?%��j�x�����5�����C�mw�hm�?JP1XK�(h�K�*O��J�l���&ᵤ����J�Fq� A�/	�~�GjA��{���z��S;`�nɖM,�O�����>�{�e�1Im N���7��^�4Ӣ��:����dX����}���5�����e��<�!L�Я��a����U:`݆��s�
�b���{Q�5����P��,u������A��r*(fI�Nb�!J�[<WQ*'����	W��R��<
{��T$��gEe1�����[m�:C�S K�f	De���w�����	'!D�4J8�v�$=���L$�k>���a�
�?с4�9�J�Q�"݆����XZK&�
�1�I��a>���:JV����I�`��Q�Xtju��[�X�g����	`ꪦ���Pܥ����^���i=5��g�~d=[����GX-7�0j����Á�W�fm�4�'m(፡g���_%|���i���J��P`�+�����6?�Ry�+5P��
~����t
�u��A��ѣI�a��{;|���o�wһ�K�<Y�\��^�Q�Ɣ~>���6Dg	�J����,R6�6�?b^-����;o]9�ԫ}2X��J4�$���y�ڊU�|�� ��L����a+�n�F�*.�-����?<� ��|��	!�u�]���|��|�e���M�;7PF6)$X�~�_ݕQ<��Nx�cb��`JΎ�1,��'��s1�+<y��T�����������G�S��>��g��I���>�K��ܲ%-������\����{p�~1Mȴ<�9���jg� �k�Glw[ h���������V�Mq�u�e�r4�����T�;m�4����K����:.��[_M(�.x�i�_i#0���ݨ��*m�y/�%��/�{y �<�����\�%��
���\N�S�V�EQ�K&���y�;+�
�ID���3uTʂ��;���j�Q�f4�K�5��w&�_'��ڝ�م�8�>3��*�t}�F_�8�	��
�x��>+���2P\��9Į\����(2�*ޔt}��x���,�g:�Ր�L��Ӹv��_N	 �JN���z���0uU��ha_�l�p69����s'�Ǿn��F��e���R�wG���$W��؂)$W��� 99Z�4`��	�z s��쿠��_��N�x8i�@��ɏ�`�4�"3E�`��J&�.�pC��_޸�6�����	��E�G �]��ܴ<?�f,����և:$$�,�)��:(�r�.�$x�с��ڞ�8����8��/V�����VFSy����v�}�/����*oһ)�$��TI�w���iFh�}d������~�8|RpØ�h����Ӊ�n�ə5��^&^8i�e)L��%�"OSo�Z�Z��bN�mY0��0��(�6a�'1s�F� P^D�m�[�ͅ��8M:�ٻnL��E`� ��o��v������ݕ��4���(]��Ʈ�"d#b���S��|@�/d����]H������U�7���V�!�Yt����̄
�a�!�~��渿F6�T��
B�R`�րɂ�� }�Q:oCD��N�zA�P��`���%����c��P�+�#�ӂ2����\������� 5�\��~��6׿���ǋ�mFcq�2�P���ȶn�k�@4��5<n�J�sW'G+:~f/����,�wM�u	N�����)�ug<ſ\>���l`�>O�9o'�Tm�;����p}W�!6T�­N�6��%A���g�qIk�����4�Y��v����9L�
��s �`�w�c.��-���3���Hl<NՂ�l߉���F��v	R2e+dGp��8�kR�&�O5���"�@1ߕ����Tb}����J[p_��S���^���QD�
w_�^^+h�T��<�U3�+3�"�w�"�j��+ (Ryo���*��pOa����[��Y��6�˘J����������2��U�뽃���\裱[]vy�Gdj����Ұ ���K4���ȫH�L:��NH������<��z
�W	)���	q[�6���z{Et,L2/�:��2�e�}��$]���8����d�b�lA�E1W`�������oQ�u��i����I�>�#��#Տ�Vo1����k�0��bH@�%��U���6o��w�ܒ�t/^�pR�M6x�6&��0���gm�Eb�L<=�X�������=F1&V��Sn̽rƅp���M>nF�L_�X&�~�����[�x����b�d�J�Q��~1v*��%�)�_����d~y��Kȕ�3��@_P�U���H�������q�s�ɒ9ۡew��-�.\�ccs�^���WY�A(�g$�a�o�N��*Dv�cY�AU6�6�K;��̒�7�|w9KA9Ɇb�bK�R�e pk��A	ǫ��Ц�#�*Te���Z1h�)�{�k��T$f����������4�!�2�&��eT��d�\a�Ъчb�W�sK�2i�!|����s����Cӡw%М��Cԋ�y�r�����Z��7\ B�~Z����X(J�=�Vm#/�Q�<p�`��ᾡ�ĺ�W��5��D��e�72�5o[��&�EL�����Y%��v�����۶.�|?J�㤕��2�1��a1����&�m8�	����P�f��z9�7�Kpq�ǹb%U	�K��Ğ`�%0
U����ݯ�����(���`T1�W	(��pcP���`h�:��/z�#d��5�/�5ĥv��?��^�$s搐�Q����F�t��!xz�����ҟ�k���6��k���_����j���q=L�i����Y��
`j��nK.�QR��PC��]��J<��zw�ÿ��O���&|�p	�.i洓M��:yn�7�`��X����)�����E��;m��
�֧�O�����L�Yޅd��
e���p��䓄�A��7w�	Ŕ����0��d�22�*���|��,�S!d�%�p�[=�hx��A��^�o�D��Of�F�M��	��� ��&��蓋3�#[�$U����Y�Xt$���o�����<�l��:��$�����^�:aJ�>Hjٯ�mű@��w!u�,s�Q/��J���V$}V��gI4q���hS'C�D#OIB�ɍ�C�-ë-�$��|�.3�O4t�lQ���9�y��o6�d�,�@x�̏sF�wHi��Y��Ń�q�����a{���N�j]hᘘD (�� � �T�Y*�{�G�Vp\C3�-o���l۽�e����w�=#O5=̌M&5ҶvfV>�~���%zF�1j��f�x�ք��5��t�֒f�����sr�;v � |�#^e�SR�wD<�R�V����9ߐ�+��i�'"u�v�;��:	�r��D�O~�v�T��$�����Y�R��>��r���r, �0�ֶ���5�)�q��yt�Q6u)u����.�����'W@*6��whbx��i}Y��Q�Nqb�?��dO<���(��X΅H�0$+J��'�+�s��N���ilo7Ac�T֖�9_jO��ƣ�����(}��� \��Mm�iaH��~�:�ݸ�����D ~�vFqנ�e>��n��ɖc�>J�f�j{��b�����!U4=n?t��8\�9b�y~1���)�)�=�u��)�p	֛��(g)_gx���l{gO�N�&p��mo��ch���}�5Q�V�R��Y'�)FY>���!p���pe!�ɳB3��o�iqa�W�5�2�&Zɇ�I|�f Y�(eE|8�rʋsmvl�l��i�x1��
ל̓9��ۆ��`�;����}�tr��&�@�k�d�FK��Jՙ�T��}Q����e淾v�LN���x�,����6�<����6}�9��f��m-s��~~��iFxF�)�Uҁ�+xx ���Hc,��Syrz?A:�����j[�s#^���K8l>t���F{��)(!���k:@#�c.��3�8e�ߡN�跊#+h�%' p���{֤�b؀Gw�� g},��Aݸ%���u}`������Vx��H��b��7�N#/ZM���E�6.�)��Ț$`��5uJ�A�Y/�Vaw�K�%(�����y���e���C9�>>&*x_�	�?�v�$�[���>ɟ�,��d�%�,"t���z~��ҋ-C�D��{�ᡃbd֭�)�oFc1� �<"}P�j���}��l�=$�0�Y�\���bt��-�6�H�'�/N�0�����j�悠Ȳ�s� ���j����U���;r�i>*������aG�E,O뱨�C� �\U7�E�@<�R̪H:g��Db"�w1c�4��'���pE�1��!j�X83���F�*<��|��� :�Cn�I�%�g
�۪�g�����5�6I��� ûQzsE��^��O�Ji+۬\G���E��6�`12ʩ@^j�<��[�t/�\9������N�.D���X��ETXH��
���Јg�?�͘{�=V ��[��Wo�yT~��9���)��"�3�٘���|���\(d$3x�[��C�݁�WZ�6���e��#j�@�
�տz�*���c�4�_����=ʵd���a��9V�{j{���z8��W��1�ҼX�r�O'}��&�]���������� �2�>�����7�}f��u5A�[S[$��l���ސRdG�.�hg�P�/������p���H@�����+�*UpzW�7�Zs�Sk�	��m�;��I"����I��WnLŬ�P�������+Z��kwD�ʇ`d�E1�\-uѽ8!�{�!g Gv������U)�Zi�ȻBw#���w�����������K~	a�}=��ͮ�T��s�6v=�;�`�z��b.>�D�B��MD��3�N_�N�}�oƸ��#���O��0�Qo�����1�<������$Q1V���˅�Ь	�v�O��q`�[m��6����i��Nי$)߁���	���EO��/�,}���;屇7�s�{	/Zs2⯤32{f�e��w縔���j���%�JW�B}��8��7�`��νD�n-���C"��zF'������Č�h��׺�{#ȯ��I�&�P�(YI�)$���:w��t$�C����=�eX'����j�]���\�1PB���g���+���l� �7�A�Rǝ��T��v�"7}ŷ�r,Puk/���	U瀙�����*�:����8�B���tz�1�ތj��x:�6�7?�qya�,~���V�?MɶZN>l�S*&����u�O�6�pMw:�na:�g=4O�"xGp��G]Ģ��BG��ΥAS��9�J�6�fۚ����8�e���'��Ț��*��D˃��&�0��V��8G�*ĵ��A�%�`
�޲aE62�VA�j�K���H���Н$�S�s� w[G�T)KҸ�2"�F��N��;�9))�+�^��SVTo�Ba��M�� n�i�q�+j�П`����=W�C�,�,I��K�w�"!6�:�v=��<��8\��:�2�Ύ����	��91:o�`ч�y��.�
���w��������H��癠z�3􅘏[�g��[����X{�5�qnMo$U�!徠��`��	s,��W���)L%� ]!�h���L���Lf϶���6�+��`f�8OެU#���i?Vk���Pc������N׷�Xا�C;H����B@,�/?v�^��F����<D|*E��`;��K8�zqs�� ��@�ykhx[�5Z2�xosʚlv�8�~7���a�0�(zvXDg�b(�4����X����fP@G�1$	�e��/ӯ@Iȍ�z�@/��#{�	A@'�^.�Qm��� ?� ��3YY{=�[}�9@�w�%�y����>#oI�2�6�0��0��l:v�_S��Z �qE�@]��f�Ͼl{tuY�K�ҭHHt���Fr��#D�c��ӍvlO�>�A��7&n���n���^x�����XP��WH��E�;��I���hl�s����0"�S$faB��f^��0�R)�2w������ԫ��h䯉zd0fg
!�Ƈ��@��
��D|��!����� r��}X7�!�����ր��)6p�OM���΅�d������?�@b��X.EI��W����tre�	oI�>�-�R���=vfe��vA�\`�p��ɤ���~��j%���Z��<��_�m5)@N����l��t��#�hf���r?R}�"���fW��Q<�.���>�5(D^���h����m07��(w_���S����$���%�n�^�+i|8��$��*��I2h� ݂.��z��/FmQֱ5��.�QL��� �����x����=;�a��H�vM��6W(��������t�w�\TI����˙�I��
)R�c?�&0���Ecr��s�@�)�������l�P��%i�'�9�;A��J\҆;�yEk�ﬓ��~�M�Po��1
�Z\GB�m���n�5G�$�
�b���w' ��	�ϳ�[Q�˒�q.��,�S����X,_dl�����l��[	�}h�e3�k%����[
��L�m
[�%R�㾊ob�7W^"�T�z�|�������R��<#���g�i�1Xuc�=E������z{�����_
�qٕ\����U������ӝ$���(U^B��5��y�sk�Fr��EySȈ�tɊ�������ܵ�rI�X��c8��B X�;�da09F�!s�m~��,�ZdvqI%�����S�<M*����O�8Jl�cnhG}u�Wi}��C�(�	dw�&/-�x�L-E�I����Q����%9Z(]�*�'w�M����#ԯϭ��.��	��4g���u4���7B�U0"h����Q��A��i��GG�öVce���er����Y��M5���X`ܩy�x�A�d]����a#�6�*����,�Y��b1,9Us<,9[U����q?��cu���^����.���� �g������oʃ�-�X��V�-i�T�و�adPg;�2�MvFRsc&^[6�:6˧�ug�j��0Aæ	}�MGGk�Y�,S#T�+�W ��6��#G��m �W�2�-���?BM~}d��Ѭ��*u��Ԓ�#���ճ�{���6���Ǥ�K7��KB��J�(��-V�mbX$"���$!�dRR�� �8_�1m'N���㶋� B�&@��i���T2:�Wh��$}�z܇�uwױ?���nd��Q�?��� ��D3�G��&8��^Y'��:Hֵ����Qcm��d�ͩ�eͶvj��-3��)�}���'D��J�qĸ8��c�3/Lh��|6��� �Uh���yw�����v�HSzzp,��#���ʌ��VG�.Ρ�h�'=�UjR�x�����`�g���=�5a�{� "��$�	�]�)Qbv�eK���Վ�������!,7����+(�/K�Z>7��	����m�aklJd*�Ӎ.��7�qEY|N.�r`*�b[��
CKFyj:Ŕ��`H6&��]�D�b^{�Є7����nF!�|X����u�2��x]B�3��O����A���Z�螫@���������JV��1:�T1?@ȼ�E	��Y:ȹG1{�y=�3�,���Vz��?��s��GJ�;��% �:�آ!Y�#�IZ�d6�z��Mr�B�2Ș��N�`�P�i��%)��fԛ�\5�E�%P
|��_ῄx0�ș�;N�!tG��5�G$.e}�Sؿ����;)�������ڮ'�yO+���~���:���i���܈|Q�Oa�+2e�CFVE��"&�/�� �(��̓�p@¬��Ǌ��)˳2��4ю>�>��	A�����'#��M"��_�>yR�I�w�r�s)b����74aR��M�� ��� pn.�OAh��S=*3���3^vǱl6#�t����!����/s�"�	CЯ*���-� �Ub�m�֑������A�"d��x�T���h�M�*�sR����n�+pp@�L�G/#f[46�_ې7�;�ZߌimBqZ����4�M1��B�
Kk��W<��!v8�K�SP�2	��}��~���F���C#2��d�~A�e �ɂ$�	FZ���إ��24"����A2`Rqo������:h9�(n����Ï:�M�F�i�,�,�+V}m-N�u�@צ�5���_'����p. 8	A� @ę��on����h������q$v�e$bU;��KvP����Š�#�� ��D`;}���虵�Y	'ڌ�����P��;��2�_�Pe�NJ�QW��0�"�/�k�.���/z���}|m����iE6P�ԗ��hQ�v�f�C�n�g��>����;<CI�i��3�1�x��k�!�F�3v�[Ѣ�i>ckO��&����T]��!g���4i��C�D����k&3?s�Y'�Q,�dZ�՞Ɉu���xM��Q9t!
�.�����, �U��$?|�Tb������'ab��98�+��UcV(��k:x��~]�W(���`)�W���	�tL>��X�X���*�H�)��F������RWK$�>h��v����z)HRR�ᾟ�	`F��K�pY��	�v;�[֬3>�O,�� �*&�x���g�k�8P%���_�� ��R���*3�qS$ף�XD)?�I�8���a�KY��H��O�Q��0�V�'�*�?�����=[{�H��aAU��H��PD�J!]��D�����q&�?/8!�Kɑmyo�dh��j��h�]��Ps{���;Sl�@�_�2y��
��3�������i���Q�yK��⽡�sixk;�w0��^��b��ly��X�9i}�7�t�hR�����W/""L*�ܲw�6�R�:xg|q0[~jǵ�zˎ�̟S��9؟ʋ�n�Vج����ǜ!vPo��$g 1[[�wD��&㖜���r(ʆsW2[�����Zj	�c�n�E��������BY��#/垑F�"l��=�(�*:�H�f�U��0�\��Ǘj8�͘R��0�������2�UG��<���i<��tj<b���+��e�ԠS����/#�.��pO��9Wd��jF� �Pa����!GbO&.�=�ޮG��c)�R�u��<��MJdpz��4�.t�8�)��Q���c�CԆ�,E,�Z/�^T���Y-1�
ڳ"Ĳb�N1"����s�h����3-�a@�&�2����x�sq��
�
�N`����Òu��^���l�'ݖ�B,�x���k�_(@sV�c<2ӂ/�{��%���#��X�:TL�M�x!���X�^���3�p�f)����`-�#��%Th9��P�)�Ec��	z�8]��Y$�ux`��l7�DpPug�^�?��+Bl�\���h�4~]�s�0X�i�_C��t��f=[�^Ĥ��9����J��<CN9M����%��T^�Y��?˩R��``�/�m����R��7�H��.h�BK��;�MOv�h�����le��	�����ץ���<4�&T�QD�3�2��+����D�ې��R90@���]�]��:��hIѰ�T%&j��،�W���y�O�O�W����KH�4٠c�񙞭�d�?��@&#_�Q�cmt&`*,�/CYfF�� �j;����.LT��U�����Ct�UЀz,\�+P0�����Iz��#�ĝ���`�B��&�,�ON);+��`K�Z�&L�/��83�P�~���B20X��KKV��V�Eaz6�m�Q$��
��������R���.�h��U���r ���/���N�w����#��+�ky|We�s��eV�"�a�Z�J�� �,�T�,iC1�]����4ԣh$�.��*J�E֖�\�.�����ƣp��X�|�Q6A6��g�M��e^��
E �?#�Q��0�Ң��m��eb}��������F8ʕ�n��fY�$��;4�X�-66���]4��9:TL
�t�������h+!`V��r3
��33݂�2%��s����-�5ڛY�	�X�"jdh�,�!���=�%!5��t��u�D�($,]�/�bBZ
�u�D?D�M�6�6,PM.5:�W��*��<�,:a�"��P�$%�	|�-�Ϋ;h�w�����I��F���o�&���9�0�<�)o�&�-
�\K���i���*��؊��ibL� Ƣy�q�Č���¦z��5�����%�e�h E:�t�s��5p䪣f�(���^ t-�ɏ��;�g|����Z:�)�s�d�"��Ӷ3Q�Q��ǥRݔ����EXXu�i��A�L�}L.�d��~�u����l?Pk)��/������c �T}\{}�j~�u~�?͚%���Ϙ>#c����/Ȍ�_�ޠ�GS%N4�[�����8�f�L#ȝŪ��(T�=S�6M�Zmg��]%=�Fs����I�a��T��N�k�(p��zB��c;�*q6�k��߯
����'wE��^�`���zH-7TB���p�����}���&�[
[�R2˹�[��d��a��*+I�g��@�齾mI���C���ŵ��w�G��Y�������ZF�mehӾt����d'x4�m�� ��"�|%�z~QF�-$����70��@'K�K[��m���៯0�:�������G=���b�a\�������T��3
)yũ$�^���]U:\.�P��~��&�BM��L���ܦՑ���.�`0�b�X`lD�|��RZ�r�������
�X�#�[����e�� ��zNc�C��ѤvKQ�r}��ˢo��I��Nze6�*��^�NU��in*޲�p���Þ��HԨ��qB�PM�gg�+o΁����׭kV���Ӥ�;���R��B[A=�l���]�/xM܉tq���<l�$𗓖n:����APJS]`S(C��W���(`�bA�P�kPj �,�ᴗ�O�9����M N19􅴀���C=������]MZ��������?.vy���]�w�>������>hOB���ʐ�{*5�^���"�s��fsvާZ�\,�*]����(١�2R�����
�+�i�ʲ�Q�lu޲���5Q�j�u9"7W^��9�!)���>����x�/dE��<d��u����6{�ЕTFx�2��x��{v�v؝�L�0n��Q��K�X�\GWƎ�-�Fy�U�ʹש���"[�=͒\��m-��-�-����+�ҔEQ�������2�/�Ԋ�����V� T�?AS��1����JrZ.��
�Vz�m-�Z�i;����l����|�	�P�I�?�(��wO�f�'��u�9.��\!��]u�����%˻��-r:�sw��B�2E!J�f�j�6d�kYr�{|&졕��趿:����LQFkX�W�s���-j�Jz����]4�P���P%RaQ�_�%�j�sPɇ2�{՘T�3�0�"ڲ:��=�MIL(��H�^M��b
� j�W_��?�\'%{n�8a�^���׶�OD;�v��F.}C�Őa������ ����rzVp���_�Ȳ�lS�
%�HU�d<�`}�)T��(܂b��)���/�A�U�S�	�IhE��<��
j%U�8�f%w��;6���V�Y�� ʺH~�?^0�Sy�?��{�:@�3I���zg�ڒ�9�Rz�)9�<n���.l�B�q�H���l�:��mf7͝MZ=�A5#ؕ�|6$�,�=3�Gk�V@ݼR��B��E���؍;J+���iA�ƨ�H���*���N׭!/�Swd�<�}��@��wď�9���1)��RL����a-���pCz 0\��0!��p>g��\w�)���P�Y���p�m��7ti��<B�X��\�.�Y��lT�,�p��%��ƹ|01?�ݗ��-B:�Kwc/e�Ya��N?0<]��� Դ�w�*�ٌ�B�QфfzT����I���s��)n����z���@�IN��lƵa���J�#�}ؤ���v}�3��	/�&-���b�<��7�'@�L_�z#/-��?a,� l$ͮ �n�b��S�V��jQ���0�V��ɉl,��S6����{����N�� PL@�w7����t��9���-�7a5l��X�pWs:��f�EG�ȁ���M��ت�'�qP��]�`-��� 5%F}��2&Jk���p����f�
G��ZX��t_Hs��g|�v�N1���j�g�"�Z.��JW	��y�ڤ�\}����CS_9WwVu�u��tJ��!���`o�\��nJ�s���(9wk,|���?KdN7�_E�/�D:V�#g�hŤ7��^�V��=9m�~d�m%�hn�;�R_yo9�ƨ�8�dD#����<�C*q�bm���u������p�/�.P�}�N<�uB�����U�6m�-�L�癆�s�|�����9���B�qyLm�w�QC���;�z+�Z0"X�>q�(z���
��h�2`!zo�H^<Ϋ첩
��a���^�D��N�I{��@j��?��LN��9�f2��芊+U�U%�]��ѡ`���<2"}�/y�mvH,lu3��Cu�k�/9�o,:���(7
�պo&���b���c�A��}Эuo����5�
5$>�6x�k��5Є��z|՞/z��/x~ML�Z���/�OԞ���!.�� +�Æ?g�����W�{����D�����
G��+\>�3�Gp���f�=Fp6L���B��N
٩2�ڣz?��Z4�R:<-�q�قs��"2Ҵ'��VY�>��T1�fUlFr�+��b�o��P�D)MVq�K#�s���:�|�&�̓����-�+��Zv����3�t��[�+[I�x�{�>L��ע�t�]l1ӟC+O��sMƄ'��]���?��ֱU�;��k�ܖ�/l^�=�Қs�U�w��D05�	r��5t��xNr�i@��j	.��fP�橁�Y�v��C���;�i$x���F�h��x��4�/7��iWk�b�{��6�����jG~��Y����?N�D�P_�V�����@�u��<�21�!���Iͻ��;w���#�-�6�V�DH+uR�SQ�:� f�܁j�yI7���#�ަ��N���Z`<�xC��2{�K$�r) jl'>T�L�L,,�Ih�a`�|�.aR���0�I��4
�������~��ǃ6��~����9��k�z��z���A)B�v|�\���5}�i]uk��#��%^Bhu����_��"M�\-�Z�`{�7�6)E��B���F���t���1�'?|���VMD�qE���;C����r�i��T���A�.�Q�V���E��$u8c�@Ki��\ա��s��3�s1&(j���zJC'�S#e�h��LxK���c����+}��h�$i��A:#~}W�ϰ�m����I;J�����3)�D������ ���2Y�v�@2��"I-x_??W\���ko�}^0`ViJ�20πK�1�Ϸ�r�:*��N�?*S�L�}#��n�zs�j�PtNN�z��y��(�$���m(T���J�[���w��_2׋�|�)�c��Y#����v���`�����UɄ=�,�*ټ��Κj��H�
�E�byBb5L� �d��UCTN�X�k�j���]
��u�j���@I��GH�Gx�2�`ǋg˄��⁜1��L0��+cQ��p����Z��@:*#�m#�Ի�_�?9wK�v۽l]��9��s�����{Lzǜq	{4GJ���8�+�0T����}�[����V��(��x-4*r/�c�,�)O�gu�d��9�$�rX}�.j ���rwxn�_6�XӰQ�5������6@u�'x����Zy%aK���q1R;�Fg�7�~xH�*A��H�1�95+X�e]��"�'7^L��^�}���>��{|��*�C�zMNngdFyC���n���%p�d�@�#����d��r���ȿ_���'76����f���b�i5��+�LTs��}�ʑ����������E���b�0���0�K�{�>`q�Y����A��U�������ok�VI˅Z�����vu�ÿ�͜�t��1�̃y����,Y���0.DUo67R�ej�}*1g&}��8�}]���~��=��y��ZKWȩHK�_���X�t[|ѳF1L8��|�|7�@S׃m�xpхE=�>�Ed�L1�ͨ �+�"
�et�� �� >������s�9�|�B�+mi��G\�S<v�A�r��C����l�<�j�j����CX���&S�K������qN�
� [�,B`�ε�m����Å���c�m�5�D_Ѩ�G��x�6���RnU���u�'�������zJJ.;�餅��~|����E
b\��RA�]��u칊���֞�g1���y�Sf�Xq	��o��X����+#�5�q6�=��Q�V0�&+��f<�~����hx3s��c��/�� �<?���5۟���'Q��H'ʉ8��+�vj5Ј2�}��M�� �qU��%��|�8b6�-v0�N�n�����r�GG�%a�
��,Q�y�tf���L�BdAQ�)]��2�����a��@(r�&]2���)2���f�m9f2���ڈ>eݗ��(��CA��r�7���춏����*�hy���$K\�R��SaY>��C����J���}��3����R��/K'A�<#T-أc������2��5��0�,VpzW��u'��u_5T���` m$am��)�c���=��gt�P.��aп ��A�Q�)G95��w����D�3��S� �����BM���n5���H�𥳎AC��ߝ�F�����m!k�p�v*8J2�I'@(k[���H@���E�[R]���T��	�"1��1��+'�N����X:��5�Β��z1"��l[�X����t�L�́��l	�҄6|��������F5i"} �p����<t9��\z{\g�l���.R�kRѸ�c?]���]]�Y�ZY�Ͼg0<�9�H���_�԰JJN�ݷ6Y�\_p�c{�x<W=a:�5�4���rB����ͺZ�r>�N@g�>�6H��1�Ժ�Q���!�SmD1
w����+�ę>��-��"ov�W�9�K�������h�xq�r��s�5�*m� �ϊǛw����O������m���.�@y����f]���~L�����1�ƌaQT�R.�5D����^|,Р�=�r&�E��6$�h��0�lq�>7<�W�!�:�����0�?���.Ppl/�W]���`�¹b.|&sdĊ�}����lme��`���@��I�QŢ�G�S~!�+E9�`i�R�l��_1���L�|������Iͮ� ��1B\�1v
ܮ�po_�&9t*GR#5�]p
;�䮏f���v�$��GA1e�b�(�Wv}M?0��@�E���I�+��E�Iŷs*����=ƒ�e���4���)z;mZl���5��~�%�L�aH
C+U�K��b��=����Fk�s�/j�T�f;c=䌫�X7
F��W���nT�L�8�ʰS����1��B�E����b��}�uޕ @^��51J͞�֌#1�|0��E6�&ߓ47���wr9-fD"_���sh4Oٶ�݈�ܞ�?��߮]�1�o�9L���oU���,:�eid˩��������e�a��Z�����M;��A��q����W� �_Ӂ<�K9�L¿e���**�7�v�!�s�X�=�h�������@��ψ���w�(>�_�$GR�zKS~�L�Z����M*��$�S�K<�� ��%����}n#y4��ź��9/�8.v��ǳ�}�����D�P���c��`��B�k$f�p��v����:M����n5 %B!�l��g�c���4F��Il�&Aq�br?~��>�C�� �����|!Cb"d)�a9{Hs匓�(� �Ce�^!�Lw(9��з�����L����yT:U~�ƿ���V/��U�T��X�b!�G���]�23�2�� �1Rb�u?�`�t1_Fd�����F6����$���@KsP��'!g��蘩������̲%yDwǚ����hN�c����zG�E��5l�2�^�J�1�ډ*�?Yo�"B��
K��vySF����=~t�P�u\�M�0+ӡ�~�d�{�_%<k�
�Z��oa��mF�� ��%��$(pOA�k�(�>vSs#P�_b�){��{'�}>p�=�m��2�I��$d�1�Z�I�l��H�%�L���JC�k#���֏a�,�e�-�++�����$.��(�QJ��׷��u����7�����#̦��FH:|�FY���Q�#SN��'{|���+*���eBB\r�q�"�\�+�04{��k��@(\�ׁ}�ioQ,�������Kc�A����V�(��M*��Ƅ��C!e!A�;�d}�O��{IW/��3݄ۺ�f��}�,�b����C]�&�%ҟh���������	�+|<)��0��s�P;���-����#K҈�Ζ�;҉=�_��T4����1�w'1��ˌbC?;��ӵrb$aTξ]��|&�|6RƲ�7H�7�K{{�w�HE?��-[��lP�Ȕ�o�_+̋��ȥJrp,�a^�`��g1�6�U|�s���3��M��k��	~���ϓS3�L`/3���l���H�x��'�n�\a�����x��Rb��a�h��� ��wK�O⃆��[?C���9�@Iro����V��֌T���U�Z���lL�+���-�Zd+�1�c������p=��4@-�{��κ)��_Jb?���N�ݕܔv�N̎<]@-�v ��j�,0o���լ�۠R��}�s��Y�o�����f�ƭ�F�
	�_S`U�Q߽Ų�22����|���F�S��	<b��Y���5 �S��7�ؑ���Q��[ ���<Fu5#���7�5&VO24��]�Yn�}]a����j��-R�pmR��M�U���CU�����xͭ�B�[�#�S����O�+L"���@�)u�۪�o!�� N�P�VB�bTD�����w��|rHU����'8J��s-�@���ذU�h��knw6�q����OP:m��A�s�;�������5����8mbq	��y>�D���~�"j
w��l�I'={�Xq��_xPR�ZC,˃i2��$�+Β�g�ȍ�Q�mٍ�\J�iVy�b��,-����nd�����Z8���^��>�S��j��ʼ!ֹZ\�O1`��8���Z��d@R$e����T/��u[`?�z+D���?��tTP���sT.ș�a��}uHG�3Bx>8��K4(D�D�'�oM���}����n�v\�9��sB��E�"/���ժ�?d�3a*�RzVM+
>ݢ�v�%��9_�>���(Z�3�|F7۶��Ƨ��o�uH{~��%��!��@ǂ���ɥ��������c��mߺ�g鳵�~�J�u�C���h�
j6.5���a��Ě��E+G��a1C���xd��$���ѺZ0�$G�Wj������ ��T���vQ_���Y��T�7��)�Lx T鑋$3�d"�ڻ]s=s����I�h��*�<;2S3%��c8�9��^�[�Oi�]����0�U���I��&#VL�6cxq@y�((��x��!Yy5QZ�����z�,'°���"�7�[�$��`�3�QGAQ+�~c<[hl�����Ŷ���<�$�D�x�����G~����v�G�7�E�|��ʐיZ?���xvԵ+��+ b�@#͒�+��L��w�����90����:��;�IN*;�����rLU5,��||w����?��=F�-F��������ΕT#��Ԯ��&�^��$}�u��ډi��5���W�Y��+cj��ШD�I�w�Ԩ�w!� �ttj�o�;��Ck%�l4\���@-:[�Z~�$ju�������������`�<߶�h¥=�eV�6MQ��c-Ex�	�|�]]R�i�+�'PI�IS�`?���F9���\���Z�k1��\�z�oL�emV�2����Īp��H���o������>�sV=\��Ӊ2�h��M۫��7���4l����ы�[���C�1#)�v�i)O���WƋ����,��Щ4��\�H��˅9]����p�7���J��q:�;D�5*���L�N(��#����#�`��xlD�$�2*:�������t���I��wH���]0�W=�y�I���HR�%���e�'TE���p������A�.�����(�B(�w=�^��}2�T��U���D9��_��
_�)D���S��_�i7���5��K��	�1ӹp16!d��Q��sv[FR;uM�hԭ��X��G1�d�IA~���E���<�֯'�WipB,�q����VnGl!'vXt�1gPZz���u�q��	�A�_-2/�� x[�`��h�ƚ����rmN�;S�v#��i��Û�0�b<���n�)+��#�aKn���?II\�ۧZǷ�5"���h���r����]\��89��B��)��l(<:�^x�N�*>�ڈ%�����ɓ�pC���ePT��6f�h}�#���i�X_[NS��YJ�!�5��57[];8���)+����?�ޕhx��m�I��.S�-=��I����J9,S�����O�(�y;�����"��da4�&�����se^M�5�mA�dm"�|^���J��|��tJ�W��}'�����A���H�C�����%c��J�a�����������`�9�537B�i���u���$�p��j���A9�R�I(�ǂQ��lR���bȅ��^�W�	1u�΃�y�!;t9rv�P��u	��kf/=Y��τ�Z��&9f~lh [� �!e=�ʂ(�iB��d+��� �9�>�.a�W���Z&�<�d4�`��#��w��x�����P$oKϭ�DS>�_�����4�m��F2�k>!|�p����rfU�ˈ6�PL��I� �a���'��F�N	.i�Yg����N�&���8�X���0�e01�vYY�0CZV�Vh�-
�y����~�r������q���k=�U[>��b�w'�qy�p�" ��
,U�^�-ӑu���ɧ��N�ɞa��4�ۖ�����(g���T��C�$�л�gn�m��~��#����n�fb��쿐�	�V w�!�U�Z�%ԣ�j����VW�t��+�7ɤ��(v��al���a��I ��mh$��V�q���)(5���lb�maiuGI�����=re��_^� ��Lp�1nŽ�2���ﲩҠ���3-����8�]�����M�( ���C=������?-I՜t�V���ok;�Q�O粩ӇgD�E�~"%��t�{�Y�P�4B����ǯ�!9���v[��	L��t�Tc�_-d�R���:�P�xa�W��*9�0s�1����K�]��T���E��5���A+�im-R��V��	T��u����u��0g�c�V������1zo���a,9���nN}::� ~;A+���(x�k��q����/��d�9���B$��ֶU��U�V�ǃ�{�2C����\鬹\.Mc7sO3�؁T�1�&f�N��ל��ʥ���/��`�$d�3q�6�	\>�hv&0�d>��-��֡�0�к!V�;�M�!~�*��y�.H"�qj#�;�f�tZ�� �.��u��?=�<���$��jɁZ��H�P���^Ǹ�Vy��`��P�<J�H���$��|͕orP��N���<�h��т����Y�0�=ʅ[�eN]ߔ�-�3 [�{c����P���r� ��˻�YY�l��֠�G�M�4֬b��bz���F�H|-�(R=C��K�2a���9�ݺ$@D���0O�IB���P�ja�Rv�\�7����%�J��\�m�T�T:�(��Xa(��S���p�`绋C�Sٛ����}�'��[*ޛ$}�?65jU�?\>�Z
����A6�hQq�iEJ�Jvfs\_5��*��ǆ�Θx'�C��r���@$u��m�N��
���,>�S\����xxķ��ܖ��b���+�Y�@6��;��� ��[#����>�
e������.��f�N�@�Y�s��� 2rؘ�>�%�]ܼ���h!þ��L����p��c�@���	1��
Te�M����(�h$�m���X=�S��xh�nYA��2v.�{E1 #9�����}2$|�ԕ/,[�5���IOV�3Y�S�p�JQ�5�\N���ڳGQ�� |xCت�����&����J��Њ� ��S��h�ϥ�4<)4�N�Z!��z@�E2��ٴ)�X��$M����߁��8���1����a"V�����3�������9�S�f�Z@sڽ�P*LOO�Ѫ(.#�*�ڰ�S�c��Q���`�L��"lr�g��>H��s*J2ޑN�%^�tLȋ�B(F���E� �Ф[�~i�n_A� .DDJ�d�H1����q��^[�ˉOB���q�S:' zi��:Y�'�ߏOFp �&7���w���h)w=Txc�45֗�=(a��B����(f�Cj�V��k�l�:Q���0Ixֲē�(	k��%��E�$�|��Z����0a
�*����@9ޣ��Fd��؂���o�̃��cJ|*-��4�	1�-
[��%Z+\1�&�WqVn���<�K5߀�/�q�Y��dQm��P���*�����z����J��B;������zu�?�BP�K�^�8ro��cх/��h�O�{Qn�a���|��0�IQi���u oE�B�J����(.UCN�}��Z~?��e44m�`p����ti��*�X`���
����3�ʌ 
��m�6p/}W�3Wޔ�����	�*A�yj˺��ۣg��,C�m%+\;n�+ZW��=�R�-���8�A���|�<L�ŔGY�1*�k�㥧��8?���{�M�*�*����F�:u�E ���uyr��:F:�(�����Ʉ�{G�X��$�/���ϣ�܈��J��qb@5MC�ܿhs��X��ӟ(���	{	��Č��R���V|�&�u[�Y�ӡ�.��{I6e!����E��@�z'i���DT�O���9^t���A&�Cm�n�:hyX X�s�=��Iy_+��4f���i+�`��OrT˛n�l�`� R"Y�"2����it��y� �R��([����q��@X���M�qv	b0��i�ɟ��MJ�A�	�<���7i���)r�}���d�S��\Cy2$6@5I'�!p)ߧ@�W�'2���Y_X	K(PZ��,�Z�U-I��+���_H~h��@8�O��.y���|=4�CB^&o&$�0�QƷ������R*5��2�6����2S|㏘wH'��4Ri�Du�I���]������S(����)�Y}�L�;ja)w~<P]t�QC������Y����&?�T��9����o���&h��V�e;���A!u��-�:��2���V�*�ʦۅ��%�5Aw�Bd*�&p�)��8V+�?'e�.N��r�Qc1�K�P\T�X S��Ut��j㨂��j� �jV�>�*�?���Dc��MeX���g%PS���R�d, ��9���)�GS�e*��L�uK%�+
�K�$�s�'.�K3�xk(s	���}(��lQ���ü��sǦ"tԟ̵@����t�.|��>�����Ʌ�K`Gr�<��n���l<�*�;�~��|����G���x��b�{���m2���?�����%Aǲ��1<ƪ��m3���>�<x�g4U撏"����̺��^��L�!��P�K���'d�#��_�<��X�i:�ҕU�����*C7h�����}$�����i|>[�vDν�����խ�>Lw1�V��	¼9idt�����u_�hp����J��r~���$�������HKJpEE���5�߲b��K�]ѷ��)��k��Bm�0�xph�Sv���
&1�I�'^!3�3+���r#}l}ߊ�Wb_������|e)�J�Kq���:-A%ɾ6eu���A�_�/�����9���R{n�G)�V^�Q2�[��_��WE����Z�,�y_��:�܁�se��8	�Guڻ�03��^� m��{η|��d��`�2��=[�VA�q~v�{�0چ��F��r�é �2�Z��ʞ�b�Af�ʳ�Nх�U��= ��:�Yij=N%�Z�^w�����j����]�e$����K��b2�.Ay�<�<��		�����.�5>���_~���W��B�1�����b��=."��ц����M��Ï3����;qwBn �R�#9��y��ߦg�����`H�O��j�_`{+�Gθ�k�?�I�Z��K/?��� ���Q#��U8�/�-ъ����+��h|�T��H�|��^	�@����5�O��'!�"�?���]YbD��ڍ�5Α�o܍�6��	�3�*��6����8��q��ZU��f��Y��|E����S��]>� ~�J���E��'���S�����9PEpY>����E{��[;�	ꑿ�a���U������}�,�J�4��wS�=ɜU��h��|�#�n��e�v�zZXZ'��9��φVD^&���p��2����@$g]L	9�
�.���1��(Sf�&���UϞ�k���ط����F��*9��O�;��NAKN��onP�>�<�<��uU7u`�հ�<R��b*Y�����1�i	#M�s&M������ق�yq�7|�d9i?9��SB�L;��o��p�0j�Ҹ����̓�/�0_,y���D��T'.��r�_����I��tu	��}S��H��9șh���Q�U� F�O��g�9�+>k:ֿWϗ��<�)�o����#�%�vh+�n�=���x���?�n9�H��������m}�g�xr��Щ��x�<����ELg��󦳲F�m�v���s����^쉹� �Y�����N!��vG��(\���`+��������m���k歜c�Y��|�Þ��ȟK���B���Hˬ�.M0�B�AW�s�
��t�I��DZZ�T^V;tW�CW[� p�{<�����T��
�UP��F~����ш)�(O�{�_*ݡ�3rZ,Q	�]�ɺ��/<v��(c�l#M��!PT��v����	��1ϫY�x����GcT�.��e/�z7	��; ӭ�֙��C�%��+;3e!�.���I�(Bb��:襛��#/Ƹ��x��5��
���9�hG���9u�������M��J�
��r�Hi�Jw#�u�r5f&t,�$�����)V�!�p��P���,���K���*��#��	�ϥ	�&��Ԙ��s�!}��E�I��v�ˌH�;F�����e���#��bw���j~��(s�ꤶ���|Ը����P͡���V�����U�_��2�k{^pD�Uh:����IHf�")1X�hp�lLU��`o��:9A���{�T2�����xo�� ǒ1?v$`1X����A\I�8sv�U�"?Q>;��:ZQ�-�9��/V��d�j,F��~�Ǒ�p>O{D�N?5���/}�x4s�kݤa6J�0a�HD�H�`mi{�a�2#�P�N�xM�ɢCA�:���^��T<��(��'mN�+�0����J 3_,�d�O�-a �펞=h����;/�Ｘx�w�*�G6m���_�ڦK�#���/��A��M�Y?
%�l�'W�k;�b�H�}[@*��
�BDp,��ٻ��a�x���l!���E~�Ɓ����=�++4wcs3/w=���+�A�b�7q�+��류�zͱ��K����F�T���;�_�� z����u�B��>
5(@%�����7G��<2g6�vе��4��_1Q�Sr��Rh�1|[.Q����+��z�9���m�/�lu���2�L5۴j5��������R�9�һ�A�9�h�k���D�C��Fo��ʿ�����������V��+��6Ғ���x�d`�}e=���m��3(ȹ��.}+w6���O���G\«%�ÞHfK�^�����6�)�bgw�3���1�x�����m�T4�[�O�%9O����.R� �j�<�&^є3�qOU�c�'��NY+���?�mY�$�0"m(&��~��i#U��;S[��+n	����vK�����y\�ah�s�r�C)p��b��MԓfB#8���$�P��� ?k�>-��<�C����P��gl�t�9V��ir\2���m"^2	��[���bQk�������Qq8@�#�Ї�'�o<v��j�v��=LX9H\�ջ�F�yFO��U�%�d녜̡��ty�N�Y��\�ڮ���B�����)�
����h�1���<-�#WM��'�x�#���N���/�TBI���|+�NB{FNr���_r�j�$�Ԓa��6���?Jl^q�F�w�Ne�X��&����-�5�3�B,#B6���T>UdC{cB�[�V6���('��>��1��t1i�}�:J�}����͒ ��v|�Z�������'ZAx�]ӳ��p���G�n��Ʊ3�� Ë=m'c��2ߏ>�h>�)2���'Ǟ�K�u���ٲ�o�K+g]/��-˵�LU�D��Ca�B\���Q��s�=NS�$�Y�w�QA����ʡw���hX�=x�7����$��QH��5���2%!8�Hk��aN�7�G�69d����}?����]P&��6= _�ix&cQ��0W�t�W�*�7�L��(�~X0�g�I���ܿD��!O s6�`�py0ah��M��'X��sm��I��fq�3n)�w0�Gs^���r<i@��Sxa�����MFV�d��L" S��^���-p̓=p7R&�-"Ky	SI�m>eM�� �F<�	O���\ިk���U������v�K��>���sO��Y�u��$���D�g�b%7e�A�}?k��ͩ���.�#Q0��?/S�_8�.YMNIr����ODm0���+9
8i���Ƞ\N�T?$KI���-�8� �/{�o/��_���1��-��%��W6�`��ß������X�YD����S�#t�$w���
�зɕ�.��|��=E���c3 ����s)�5�H�+���A��/p�UrPr��8��O:��}M�B,9i�	v�ǉ��J+���R���hs3$_O^Q+9�啣�lqȒ�3�G��!��$���|�������)>���(��
3�`�s�p?�3�%��^!��Ѳ���Y����=�P&��ml�7�
o���Aw�Z�yUQ��u����t���遆R�ѽ��}lo�ىA^6,5>'�> Q<�n?7Y^��ꨩ���Z�����e��!��v��������T��:_IX~�f�u�Bw��h��-Bl���ќ5.@�To�/V﹒,�"���Tn�|��8r��4L�H��C�iU� �,���@k������9|t)��*�XE�H_�߉!J����{�y3|�*F���?�
t>����[ӧӹ�Gj͌��L�"�'c���LA��:cL���K��n6�WI�oO:Q�3G��<;x����i�~*T�M��:�������kȅ>X�@KB��ۤ�pqP���[h�]���N�fq�#
����d�z���˃R0�����9�R����i�:SIۆ-|��Rgɸ��K�b }�$�^����o_c�b^t� ����(��U9�K�_�	�����5폁��K�`mI�~�lI��mݎ1�>�+��{���7�#�[����)�UsMY��U�kq"�����Ac����Oq��O�a�l�xg̏[Uۑ_�)2k@v�躀������J�ܴN�8}������]Q��!�,*Fz��Y�Ǧ|���VO�@;Ɏ5��k�*����cN�D�aÁ�ϰ�5��&&h��fOg�E�����껙�a�N-/>V���+u��C���Vt��������'�MI"�e(��3rU$���uLw5�^g��^r+�G���[��V�j��Z0����!��9�,��[c�.#p��ʻΣ�����bD�
�)�D�����Ϋ�����T�]��Ib��B��Y�nd����iU��P�!9k+r��uO�WP��=�PO��ۅ��{J�?Srs5�I�(�
�Z���}D�P��8l0ՠ��e���V؅�Y_��2�o�)/n�͆̷8#�� @A]�.��s��c���K��ضd��)�������|���:� �� #%�*�s�� H�:R�%	�}fW�tpI��+���Y��ZJ�\��-�ۑ�g\��N'=O|��?��@���������:"n?^4Y��z
ݒ@��
�3lX%�VݫT��D+��u���n҆
�L�*��4Q���l����W�go��*�<���,��$}�����*���v�^�� �8|��1�G��L��`�P���rQ&��}i�9����w�fR�ݯ�Nש&�
� �V��m@[��H�9�U^��J�u�+3o��E������e�����8��'\X(�ÒɓҀo��h��nU"�<�aK�I����er�e��3�Z}Vն�s�{͉"�V���p��>��vo����hF��c�b�ǌ|�MK��E��'�HN�:��o�r����k� 0����ӄ �`�D�`��{E��U4C( ´e[�1��q�d���Y��i_��6�~�_�r�vō9�5E�ʔN���s�5���2� ݑ�!�T��6�}Ńtڷȍ����	�9����D�a�Z��/�~��p>$7ᎡܸDS�U��	��*=s�5������y/����ϔP����˖u�k�� Kqa�A�m�˧i������c���#kz����'|�q�i}*��H���d�X+�Β�� E4��V1s�6�����
��\�@鏝���Ŷ�E9�S��?�g����%k�a�%���F�Ƭ�wDx�(�6kO>�'=����-<`V0GL؝{̛�$u����H(Ʉ��Y�&V�>�d����H�T������b���N:���Z�as��{��� $�+��`9��ۖ�sn���	b�B�0�����7+�"�V;4ۣȷLc`}T���T'������Ӏ�+^P׌�U|FP�G�m��,}j^{ۓ��f�-���̃�@�$��Ձ0Q�kI�q�B�á�u^��(��v�7��H�4Ͳ��lw���"|/)
��e]^6]��x����G��l� D���h��Lu�㕴�O�#�_&G�鉼����ѝ���c�H����ȂO����
	o����w+3�mb��u�k��c�C������
��j \.t��m����̉�R]&�,ly�v;����kΠU%yz��Mt����(8����S�@Z} R��������H E@ۆT��O�H��@��i�tHZ%� U0)�PF�-F�̞O7Gp����'�pJ"FC��
�z@˴G-�wy�>?4s`������$�$\ok`��$(�/4�P87������ ��o�N�����5�Wa�q�&��em1&�m!(�;�@�<��~1^"���`��d�W/X�XɈ�0v�J��.�K�S��ga�5{JĨm*�Wb����jԗ�ؗJ���#��G8h"�M��ۆ>��E��xlI�>|<��8my�ǅNNh2aZ�R"����U�^�s��T�5��_(\�npC��@��Z,�po��W�LNO@FA>꽌x�2��+�lg��#v�og��fw]��1^ ��[��"]&��/,�|�-j%�r���/�i�5�k�2�/�-]?��Ҧ4�e��J�m��CV���BZ��@�([)�𥚤�֮��fL��E�X�G��X��.^R�ߗT'�_N��,���v����A>N�w΄(p(��̆'�>�����S��b�.������7��htΖ<�~!�^���\��J�ï㽩j�����,�D�������>0�,bc�O�|hL�4��{�>�-ɬc��f5]�Q�� U�X%��T!�t�W.��1og��(\R�K),t�!����L��u-GO���rq��/V��rs4�ӷbg��"�F˺;��}�R� ��K��~��ai@q,���Y"���p���6gF&�eY~�uh$g���#����|s���<��mnO52��#���It5�6�,�kH(�;G��m�`�EZc��<�x�\�_ˇb��"2�?�au����u����d@�/�t������y��碡w=IoZ݋��+�eޠ�a\#Ӕ?U�����g��z�����)�Q�xs(�^��K�^��(�3M'-�J��;7�)T1�QG �A�'	��${O�Y4�w#j�d3p�5rE&(�P��<�w��.9t_��	�Dk�A�+�=����@z�2�3�ˀ��	f,���{2XȔj4��`������ {̇�-���XH��)pa��J�6fj�2�p�F��4���:�Z��}+Eu-�K�2~�i'��k�c�^�������bMy-�sU�PF*p��u�i2da�c�}2?�n�ݫ�҆���n�_��e�SA����R�-�W�6�U
����񮠕+���x��7�!ŀ�K�!8h�y�C �@���Ҿ�����?��s6��a��b~a�:���n��^����8�~��O�Q' �dLv`����A�_P�l�k��g6�6���TE���p*��$���찏��$%�C��_�x����<�H"0ң:�I�X`ho��Ϸne��"�������Q�q��&�p~��k廙��H7L�E�,�z��iwS!v?-���&?��d���{����m�s�x��3.�J�x�&5#�H�_�����)^�X����-V��qt�BAQRt��iT��Y��y='^���X��~t���d�����Nz��hcnf��rj�
�����O�������=�\`$�H�Hm휥uM�Y��1L��a� �(�z���F�>R��j_��y����^���J���ԟ9]ѣ�ڥ0w��r��g�{R��i�,��`	E�_g, 3nU|؟v/�m���<i��J�h�Ђ��K_#�uH�\�d��u�������f�@�8�_�|�~�T�����/,�|�'�5G�}
<�&���Jz�dL�s��OvA�8/���џ,�V�l]��J�y�f!\e�RZ�H���n	F��v5Ջ :a-?]	s�V]zkGl��c��-g��P��2���wY�k�������-ܞ=��I�F��b�\OU��3��!��6����e�s�0��_�h=��E�����֫]b����h=
ě��1��Y�m��=Q�Mг�������`��nUg���n�"��$�VH\	僁C��Z'`YUq�ҠTr	��T/��m�.��"��O�sG�m�X������/ZPNg"La�
����|�,�l?_��$�X���N�~ג��I�a( Z�U���CU�DtF�_Q�M�S�
��_[��6AO�n�)��R�YV�NS<��M/���+�J��y��!�Uھ�5��LR��6��G�r��Ӟ��w^l�7���G6�a�O�P�0Rp!}�j=�_���{�����~҆F�ʐ��,I��!]���8����jf��Z�*i���<��YT�暒K��/Ȕ�y{Q���e-�`Cu��[��$~��� ̫7���!_���,�ZЪ���̖����Rҫ@_	����	T�
��F�e�+w)u�g+���K�z=.]"[��`�W�&�u.�b
a� j�3�!�unrQ�&���m`� �q����H�pC!7�S��b�TL}�q/����ek%�b)� hGs9�|��B��C5�l��+=�1єF����Ct0/��>�ZCJ��� �'\�1�0UVaK'�O��߰�a��?~�G���Rl�v��`҇0��Ѡ��W^{�&�7�:����1���:�Dg�Xs=�<���'ϕF�+���/@����y�}��v�M0�eS��#���ꆅ�2,�M�0�١&�A�U#�|��7e����]���J�<_CT��v��9^�>���%*�` C��.Xa�X�IEw�Y��?уU_���9�6���[��_]G<B(���va��[�ϊZ-�P�ۆ�tF¥�9�4�yB� M���S�<u�$��U�4��X�E�� �[ W�|�Tg�*�����	K-�;�R^)�H� ݛ�K�arF�Q%�S[OT<҆p��t�۠���F�����}��9���c�kQ���t�x����۟���s�^��������!5�l+m>��&� �����c�T7 I�[�����6e浶�"e�^�	7۬<r�����5���q�m��b��)��a���_P�Q�«)�`
���(�&,7�n/�*둉Q-|�j����|X����or����FX���8�}h] dJ<s)��B�Rf)� a���^-�>..�w��\ ��D|�{��`bx�.�x׺,]zr+z��KĮ�
�Vt�v�M�m��k��'�0�:2oT��Xx�Fg�����.m�6��^$�d5�WOW����<1�9���d����#M�Ϛ�g2�qi����o��xx%p}��|ԗ^aD�R}`�+-���O�?�m�Z0a��3�m`���?I[��9ʌ��	M�t	YF��'Y`��g �XT�K`��Ak�$��Jpe	_��X4\�y}���&]F۸!�&.��U���'�4=Åbԩ�m3Ǽ��~��(#)Q�ZFL�Z�6@��h��w� ���1f/�9�j8pL�� ���{�=+�$|O��6�> ���g��#�oJ-ه��jn+�= ��e����$���X�8Ew���xv������$R���sľ�O��̩�yD���3�'q�-�#�/��wP繊N��ͫ&:d'1"B�d�/:]��Nk�4���oR�)Q�K�wQ�k�{��<���%�/�^�fSeJ�~�����>���;���f��qV�-���)��H�R2�nX�������W���Tb�[��n�Α�k[Y� _ITh��9��>��$�V�p��V�d�chL��`�Ky&[�i�f3A�y�V����L>!އ刕o��&�QlSZ��:�5���p�^>�܀$��:Iʠ�ka�v>�ˇ]������k�[���s�ŗ��%8�k����A7vU������1_H�`t����c��K ����8Ȩ��k��!���������7�."�}��ֽ/�װ_Q�����jπ�ev��ht¯���ˀ��[b����l�	�������#�&0�����BX��Te��zP0P���&��{�L}TM+���b�=i�ަvV��ÝX�2?h�*�c�~ �QUt��m��1*fah_�����ae�b�E7�P�T�!Zi��{��-x�L]����$WT��J���*Gbt7�8uY���/�FZY=MϤK�~�ڧ�܍�^�)SSa^5R	}GV()�_��:��*�jX�A��~����X$Dew����e��=�ߛ�x#�)?x� �A��"7_���2~��2�`��~��GTr�2��{�^���4���&F��j�y���1L. ǆ=��P�H�+����f���O��U��2�ޭ���%Ɲ�A:��3�wR,�r�w�V���݆�����q߉E�V�ܢS�Q��V�U->�>W1�#���i�n��H~�����N��$c��GqW�(xb43<0��G�b��j��"���I��
ͮ�WCk��Up�D�S���Vy�
V�q�X�_ �NVg�`N 9����}�M�T��d���K�K{4)8���
6���g���2;�g!w�=����r'ǵ��΋��
>����%�;	��L���h�q��c(�5��s�/�,&��'�X#�4���?��d�71!���`�{��&^4h���/߸�hf����{N �H��5����;˨��n�e*M���ةj�G5��dj}n�a��͟Nqn�0c��1��a	̻���&@N�ˀ� Djw-�� ZTs�8j�｟h�|��f�f��o�)}i߰�G���~c"����ʔ3�g�cy5�k���dHHЂ���%���Y�+��<O�i���N�f]����L�ܦ�O�MT)d��[8��@*YŬ\�s���#��$��+�v���cQNQl���6@4����_��Ց ��Pz����U%�N9���W����׀F�V��p�4���߫�Q��X������q���QkE;g �x�� )�#Rs�[X刡}Olo��2u��_�Z�0���^��u���5�<s�D��<��2vuOJEz��o��`%%�B��ܟ��49����[\?�łfф�&*�`�G#�nYN�A�%�q�<y~�a+��[Ĥ�h���$B]����ds\м���w[�݀�{,��]���_ݛy�_w����j�6�f��g�����^y&�����ir`-��u������`.��aY�W|uO�O=���Q���ѝ2|��ưVd]Єsj@�hxk��`I��V�Zm����.T�.ѡ��{��"�r�!ͪk��.[�e��T�Rl�nNF��)%t���/"֝�x��`���d�{�8Y�7���$�G����J�մj*�]�?��T���YY�@\ƻe��A�x�P�-F�N@}>}.���v}O&�zdLSa�����6Dp��5M����RT2��*u���f����|?Iu_ �N'e {�ٟ���I,�6�2<�`����F�,ܝ��*2;Wm�5��ǼD�$��-½A =�q$ݎ���G��j�T��&2�C	�~�M�8��2Xű��r��Z����/�}p'0ƽ(�9�DC�� о��ڜa��L��:���V4��}:�hg��ği�=����I���0�*�֥Hp���p�����*���M�9r��%��������sQ��D&rc���C��E˽_��$'��)4�콥�F�Y����7�N7*��{=���3h�/PݴE&��~ƾ��^��c&�9����u k��.W�����ۗخR�Y��DgsϾ��[�ʘ;��R��iJ���$X��$,�hn��}�����)�+�:`yu%�C�wP}2���n�B~���}�yw~������X�;f�.j��_62�'��Gzo�:�ڶ8ۣBQ쎢�����с�����5����ڥ/b���4�x��Y���epA�l��Y6r�N
1/���:��S9d�cM� ��2����˄�z��[n0����z�,�_A}Lzh�]�����TM��w�����ydl7(�Ӻ��� ����VQ'�T)�>�n���N˺c��x��A���{M�ӂG�ԣ2~�w�f������z��xp��;v�HބAD/�4~�x�]K�ĸ��Y�`8q�u�d7�!�T}F�]H�4pI2�V�Q����8,��@�rKrt�Z9���\Ȼ���~(H7�S161-���N����95_��Uԑ�|��=�fa��^WmH�1�ۚ�?�e�D_r����^���|#c�;F����2*�u]��@2�l�U�̀�cw���>��ozr!�,Y{�fb�	�"_X=D�Ds(�Y�.�O�ྊ��k���AiO[�u@������%��������dGc��N�H�s,g|Th�$�C��U'}��-8/��+Ysd�����ؤ�p}�D, :<h:��|�ek'a�8n�1��7*O�-+�u��y�y��3%�G�"*�����q����ی�x9���EJR5�Cu��� L��Ĕ�WP_�4�̾�G��!��f:�	T��R;�Y��'B�����N
}�<�싴
�}�7�|�|
k:B��=c,�;wۭ��2اS��BU��1�o���V[\�KYGJ�~���8�kw���Q	�S|Xiq &fڄ�2Tͦ���"F�D}'ְ'�6�x�@��j9@�;��f���{i��ρ��p5萐%��Z���	�MdL��v��CJ���������y������V�8&U5IX�C��� ��QG��ζE|��5$﬙���d1�"Ã���f�.b:?E���h�F�� �ԟ7�Z`���sƽ(��iX�샌lu_�90�T�3�C�����W@�)�]�%�nVC�G%+������d���%�D�����^J��DN�=��l�:w8A3oO�R�C�wuf��Rw|��N�3�[�!�]� id�p�����?����%[s�H]����V@aH2�B�����u ��;|S�aV���Չ%�d����l3�h��Hb�_�5�!��Fcך?��m�f��:�=�gJ���G�ef�T<N�=�ٺ���f"�W q*bW2G���6~ 5�z��aEl�s����WB��:�_E5����a
�ͪ$��l.���d6�c�i<I�oPu�J��\TLV?h]T����/���?=PC8�o*������Y���8b�_�l��m&{����#5�%j�z�n�38s&wF���U$ї���Y�8�I0����:ZVoBv �lc���Μ����)��ϧ��Slz�0pQ�m˱E>��9�y%����GY)�d���xk�U��G�2֘wB���W1��&8/W}�Rb[��NX&�k�Vo|��zSG��<��!=��~��m��^�7t�pv���ͣED	=�D�,d32�݃���W^�6չ��r����3�f��8�E��Wj��hɈ��@�&noʘ�5��v���9�5z/)��\�C�P����	��7v@��>%�tm3K�5 n�ڢ��5�HZB�"y�����nF�=ẇ=�y!=t���n�-�����[i�B���-'��B��;�W�1?t/�B�;�\���?!��mz�����B�ȋ^~R"�X���$��~����jc�I�6 ����s�um�C�[� (��*�D��d\�(�����*i����ճ��o��\��܏𑆆x�,�����)��Di���-;-�<��BX�qʀ���1��y��z�J���'�}ާD�*50Zx�o8D<'6N�l��k@��,����SxP1�g��[1��a����B�"tу�\��t��bkf��笟.�����P�!ހZ�O/� i���4�
�fd���3L���������m=/U�;o�k���Qh�ހ�T���t�ϵ�g=��Z;(�?�q6����5�n�Y��Քb�{b�{}u����4�;,�8��d�����^�>'��_��t�9m��:�I���Q��%�p�p1��a"��D}{Bi�}�KSvэ����\B�z�Mu�����·��]�"�`�D�CDr��N�͚�C�W[A�{]aR:�}�n��M�Dw���"A����S݇59�s��q*:�f\F��3x[�oT&�FR��Y�P�*+��\�5��n�fa�H��0ș���%�����O�+����N*@��kA�|��c!����?��[��ڱ�:"¿��A0��1�H0W�[���
��ʲ%�Y]lo�Z6Qdc�c|�zb�J��j��Y�q(�s}{b��VB�x�M��?<�IIj��Z�sLz�����By�j*�cf ����H^QQ/��N,�6j5�m�@��J���E�ys�p��\���zؽ2��mc�(b���}�KzA�y�f�bTP���hQS�ɶ{������l�����PB_z?�v8��$��}���-�t�'���q�˙iL	�/t	q�L���ǡ���}ػh"�W=6
�b�G�oF�+Th&�&߷@o:Q=�eL��YƺH.�ŉ�c+W�g�(Sl�����S�Aw�$
ofF�rD
)V𜵾�h��� |L"xq����-�=��n��R�!w��/��J&F�y��'b"u�d����]͠u=�p�r�ЀQvz끢_4�z����_��z͋���dֻqP��<�\��_�����*�v{�fAۣ`0�>:��ڴx��"L��T�ۧ�����^�I2$���0<�V��]���h�記��B��~SH5�}����U�;ږ��` w��[�|I)�#��@��j�2�G2�Z�p�'�}����H������S�.���:��=y� ~8}D,+/� �h`���5%P�8(�`��:�am"�Ƚ��%wUEƼ�k�~��W.Z���}6��z��m����K}.��f�Pu��Y��4���ޜ0�@:��=���/bP��z�	d����݈^��4߹SM7��_��W��vЌc�~���
�j�$H�sǬ���C��Eo��^ʬ��M�K
�J�^6�B.���D�h����g�))} �@cF\�w6]E<���j��ֲaT���"+d�"b�n_Y �G]�;�◩
5����I�ZI("��)�о�?����[�\����΍|�8a:,N��K'H}U�5-��/�˨Gj@c�L��fv��g�R/)<�&wF�t!�pՖ/\�<�������5?��n�!ћ�K࠳D1��9\�_�����?M�th�W�Ս��7t�:��Kˏ	6���r�WH�O��i�s�9��0z��4�+��C!�+�V��Ԧ�
b�c�@_����9�-�_ˋ�E�ZU]S��LH�v^�H�qB��+����voљ<<��Ϟ\���U��Xw�@_��w�D��Z�>�p�k��q�y��6�����v��M+��g�^�ș�d�P��aJ�Q������཯��J���Uk���g��l},��ڇ<�1��`uX����R0��:����#H0a3vy����ܫh:/g���Q��魦*� +����]�~[܊�ϖu@��!"�$�97���h��$���Z�J>Q}�*
�������²|er�	�Tw�?�LZw^/2'���n�+M|{�h�*��@}������(6Xy���w+�Z���2Vr�vT׆��\�@Ν�;byL硃��3N���}Dʅ�K`=B$���_x�@]�q����4�҉:����ā���Ic_5�xK�͗@�FA���)x��f��t���:Q��ڣ�F�;�o�%�p����]�N4�<����E�ꯧ��U��P�TC�w572]�j��3�Q�����Z�{����C��@�AP|8�j�L�!�R�U���L�*S��Z�d RK9�d5e��F��O��ڷ�Tq�� ����`�q�-s���mXM�B�K?^�Kk���������P���x��)	�M?I4	�␗:��I8�jW뺊W���1�f}�QHy�Fۮ�=�n{1� ^C}��N!��ut�J�{-�w�	~
�E��N���������U�ؒ�i�gk�W�%�oyVqğ4�u_��X,��TQ�A(�fg�����r��2¾��n�'�����'��V-�N.�t���>xf��#$Q��z�g6�Sٙ�bs�;�O�)`��튊X���b�4��æ�\��,3��̒��Zr�	�9��>�J¥B��Sl�ߪ[��[D1N��*#^�,ڮ�Lr#7��aZY��z���tk}�f�n���>�|ߥ��H�����i�W���c��s��W�j��H��A�����˗`����궂�f�jS��u�O�C��G-�
e�U�4�C���#�-�jL|:���-�B�I˼��^#2�ժ��~��$�Q"@#����RB���D,<��﫵y$��<�?Q*�w| ;�/�hV��k
P\=�sN0��Ќ����5F� ��Z<Auc4�4M0�Ļr��~�}󯧆Ԛ=�O�:6u��p�'��}�40~�4V.��j�ǘ�t��8��?�0�F�.T�\��U�Z�k���q���t2�4��ˋ[�aC"�ӹ/r�b�I�Ӷ/R�t����] Ь�XřҮp����4�"��[Ϗ�0���;/a��dԘN�f�J���ʄ�`��yc�N����~����ߩ9��o�����!�m	 '4{�k(O)`f�jg��֏�o�>@��[^�ض��e�=p��tA���!��m�W�Y�C��w�j�T����✼_"Um6J���C���]7Ҍ�C-���73�-<����c;�86�U�'&��p�:�+���x�-5�	|B�s�4�����)(�D�ic�QSL��C24��Q��B	�Aw�IԻ��)���O%���R8q'�,�8c��@m���j��mT	����-bk22�O]r�ǭ��Tcb�!�v���t��
�"��֦*����
�����p2K  ^���Qi9��m�鎣�YT��E,�[�+?�~<W�tn�^x�WΤ���)^�����378�I�<�]�^��4ol�y���� ��ek�^A�ݯ�-��!�`��$���5�b���^T�'D�S�]��`��׸l��Y��&B��ݭ"N[���Y$����u�7���bb�5�����0S��m��-wЦ�}�,^T0��d����q~v	A�p���[U��j��l�H ��0���X��O��Tb�o��򓄜���+��Sٽd����Fr�����x5>po��MX9����Dˀ��>eBؼ�����sg�\��苼L���|j�Z�h��U<���'��W�N<v�g�Ԏ	y������o5�ԨN������o�mz�˱���( �R�I���&X�m�OC�'>���'H3]ɕA,Bl
��� s�KG�ت�R�1�1�����}&������{���R�bj�#�pʤbOVV�
ȞAf��o0Џ|�ۋ5Dv�[o�ڬUF]��ǐ�"��n�p�������E	��	��W��)�d٫>k���P�3 �V�?p �}�`TU�����b?��a'�eE�,���Vh��7S��oT��ZY��E��cF��W^ܫ�R�}ݖ��My��/W]ߨ��5^�N���xq�~k��#ߔ?D��{=	v6����� O�����X}����$�ׇ bِB�\(n9�<�9�|���M s^�K[�Q�L	�JYrl�xΙl$,�)�����\Y��;+r�j�|ѕ�I!��]X��������G<Z:vj{���0V|8�%��X�]���n�#'�9M%
���{�\ZeMo!���u�R������X4:�U�~Ӛ�K'�l�r����]9K�|����a�#k���v�S��>s#b��V�;bS��^`��0j~�N���>��o��wl�nVހO���*��QG��z4E��~n����_�r��"���,l���S=tyEuM��aR�YБ8�>v���"�Gb	`�X��9��ل�;Rn���ƚ�hq�Z�v�RW�OC�0ۙ�I�v���Ў*�L>�6�K�W���F�t���7\��$N]�'?�3W[v�4"*�{d��׻��;�q���}� � ,�6�Pq�W&��;�"���/.g��K���� �Iw�}���^�A6��.��0�����KwddŐ�)ͅێ����+�S^���IL�� =d򰙥"��td� WTo��"�wL%kU�>��`zIS�G��D�jJ�'숪H��'A��.�I3vVy8]��w�T�[�&�����ZM �Q����HP���W�0&\�[tYc�b&��F�D���e�*�"�c�ԯ��=g",�k��j�����ԕuZ���5k��`o�{+VI$�A��ixRe�lr�߈��a�����å���k���0%?|�PS�,@�_�L��'����c>1�E�C�CZ�w���F/�J�tA�ѱ�u��&h:=���pr`3ڎ���S����+ˮ���#F:թcXѾ�������m�Bm0@-Ӄ�<5�݅^L��g���j�g�'S�i^t?���3�MB���8�:�WHb��V�><U���f�[W���A5٩0�_�D�'I{�Re�vdS��8Q���"gHH�j�}A�HwKXxB�k���MS	M*�u��y��^�K�������!���t�k��ݬ�G*q���2j��:6���B�߯hj��N��>�G��0�g#0r�����^Uu��(�(l���A��!�d�D�/~��=��]2�s�s=�1n���y��4T����%� s���O�W�q����=��U�*.qp�%��R�������� ��:������b�������P&N�������^g8	2��~c�?0��q�0��֦,V�n���y�@���&��`�;8<K�t���}��Ϙ���F����	�����(Q��u@�y�}��&�ɸ̞a�Pw��qt���x2��zu�����������ˌ9pC�e6g����m{�r�1U=$���9SY���tfp6˽_g�K��$zA �C9,���A.��ꭽ%7ǧ�"��^�\���S�.�v�����֙"ڠ܀�Y�׬u��> �"l�&���?��1�X���YxEK�EeҠ�zs�Z�K"=�[W!m�8��D��;"?��҆�lҶ�O�uq'��pY[@�4�>�� ���y���ߔ�+�鋳��F^d��rqۋ�3^�Hg��a�(V߿�"� t����@���jqU���x2kD�����7͉�dI�������V�A�����\F[¸cz(,��s|K�*�-�P#���'F�pO���WV����[��z��J�`-�Ƶ፲c|�m�Ǚ���8~I��<�;:������"�l��B��������\Dىx�.�8���JTp�;�/-쾁�f}�Y���B��l"��$W����0�õ���`.�O��.ʭz��pnA<��8J�EQ�����7�s�6%=>���Z�;h$�����g���U����"5�
x�$�B���Hdt-��L)�T,|-���3�B��5�f�Q/�k	l��i�*�4-�s�-��Vȳ?� ܀b'Ә5�p�G&� �	�l���փ�Kѕ=�:w7īl�}�2_�U�6����|X\�����(_�����W�(Y�M889�6�>![����t��k�UNkD�����p����LN��b����E����3<�V
�� �	kI�d�07YcZy�0����N�q3�ԘE�u]��7��_ʺ?�2��D�J�Ru:�Gy�<C�f}�`Ri=?��+���<Z��bS�^��mu!�@��&y� {X���PҰ\��b���3�F �f)���[���iVj��Z@��T);��qy��GC�9k�Rg����C�J0Q�&��45Pd{��R@�9A&��脹��O��o�q�[>Uz�m~g��N�6~�s���S���땝��� �C�(�<�-��	fT��p���8��c An���y��Oy�P�h�G}��~��+r��ߨs�S�r�XK$�Ø�jQ���h�V��OO�kY��i�2n����>A\� ��IR��OB���F��R�)�nnGk�s��N׾����Gc��{���?~@-�3T��}8��f\+��y�7	��& �Ř� �->�R�<-�Ŧ:	/Pwש���[l��ӊ���X����+r��|�t����	��MqUS@�vo�zIؓa���|Y*-�������F�7O��x���T�dx�8z�#���)��6786Pm�w��������5(n�$��?���0�/K��:��=%t�K~����> Hƈx��I�i����T�~Y��a���X��M �3@�&��u�h��:�K��Ѓ�9R�<���٫��G���< ��C烽�y~j�&�`{a�G` <t���P�>0�� "7�:�ч׮͐�������8�.�f?9�]͸�Av6�������u�+O���Y赭�4�E��Q��@�_w���Z�a<�4LѴ^�x����v!�Oy�ƪ�/G�[S�=�џ�ll(|v��1&��2{]�4��3�EOJ�,��W3��"Ki�D��9d�/qa|?FC}R��Hd�&�D�6����\c6#Z��9)��|�$��}�M�=���M�@�P�G��)F'��f��Y��<7�lg��̥� q'N`�	0���W����(���m~)F�_Ԅ6����*G�� �2���1��>��K'����9f�[�r��\�����]�/�Pcbn�n�q{g�L�x,t�	���1�A��W�l��9l��\0����Llh����{FQHY�۬ۄ�W����noMa�xTCt�����Խ���\i��RY�%����?��tx8sQ��Q9y�(�`kw��P�1,�WJ�\���Z��]�*n�K�-lI�4L���V"=.Y�N �8�P7��QUr�K���J���ܛd{e�\B8�G�2?d$5�QNq<"�k:\)�ͬ<Iv&\�J8�y�O.E��Pޔ2�ܬL�W�xF���&�K\�(��<=e�$S�Ql�e���E�'3:.SZ��9 �x�gՐ��Ր4�@�A���2�3�7�O.E� ��e*����/�������0��)�I�),����h ],s =$��Οk���#o>P��؁���(��5h��{��Vz���Ϡ�X�:�QțFu�'���1��Ӻdg��o*���m[��W��o�oBh����ȡ��m
�����99Nx�N��:�}=�Z�����x�uc�H�����2� w��Iu�,���Y��-eR ��zu�龸^�=�����!��O��)b�+��8/���]�Ֆ�~lZWa<�1s�`��[] �(;�~����y�s
���We	�[�����%B�UPHr�'W����&)���������f%�쎪��r�G�+�+�b���J'
��q������j���ʼ8/�7@�ul�M�v�lH!Nܐ�zH���a��:��������_��*l�ӝ��~,��q���Od:B"G��{eڨg{�M���n��WQ{B[����F�`Fgߺ�u^/K�κ���L��߿�?�]A>,L�?�\p�<l�F�Y 	���3����,W�Iz�2&�\��#�2h����N���a���7�8S{0��n�Bhi��z�<%J�}�B_*ir���J
;er(�������uT�C�`� m���1��|:(�)�1�B�Qo�3�*�)gP՞���}h-��� n�ҭa$��\3�?��k$	��G@$-q�/{zwߛ�B�}�Rž��rR�3����DcHU\�a�+��fN�jK���x��#�s��k�}������lQ�{$�q�>��,)n
��E�����福?��x+�G�qm�c�!�N<G��7�fF�L�l�D��Z��??R3C�5m������-��ރmw�\f���6:��q��u�J�g?>�4�}�i�͌��l�����+�@����`cNt�}���n��.Y51+}A���.��baC���}��qZ|,��Z�>��(~��̩�9Jެ�9���@R[ޠ�	��4#�|��:��F��M��d��퓎Y�ܭd0@{}�Y>�� �r�eRj��UToh!~R���'�Ř[W��4K8�k�=/��Ȇ�U�d���_fՒ���u4�e^39�T��gA�a�_�60��] �&��G/��vK�|||9����P�>kKG$�5`�,�U�+�&�Y��fz������䬨�/�H�Z�J��p�����q0Q����`�(bЍy&�*�X�o�qО0g���d��Q���,5�'��f_�;%��lM��)n��7k^���:Vdǿ���1g� �����bf��N{��q����wc�t��F�Hl��"Ԏ`����aD'�4[����sf��ϗ'pǾC}P�R��D�m���$uE�V�?��؄}�YBV�]�l7|��w��2�U�_/ݬ(ߒwkp!:#y�6R��� !s��䉘$Y�>
��߇ߐ[�W���n�7��-	e�Yj�\���u���#1�cd&*.�������sC	pK�t��W�c�� M��栳��8�yh�3�*���\j�п�l�S�����Kw���-T�����Jd�jį��y�J�~�6�j���~�F�/�J��@ᤋ�R��_%S�/���5j��CY~Kg���Ka2Ͱ�㥼ݒy�u?K�6>w���`�͏�u�{__��n���l�_=2ς�<��+�4>���?���Wꓱ9�&��n����;�$�e�?X93E3e,� �j/�hf���Z�K�Z�����}�[�Ռ������*qKM���V��2��pԈ]�jz��|��'w
#���9��"��$��#���
.R�K�3�H�C+]���D��n�"]��ǂk�]J���qM{������,LJ# ���"���Z��|$��(_9��6�dNk��`�N�����\n���8�b�Q�\lx+�,ܾ?<:�v_�@�6�������a�L(N�����Ҙ���9�X>$�D�-�p�ߪ�����ns���)���D0���i�T��8S�}�R�ۤ{��+6K3? V(��;�����|� i��$a�o�Il���x#(���(!�<�?�v޿�$�t,��Kk�,+6�j�|�V��Nj�ܞ���5o@�ЯW���-��%S�6�h�"�4*��r]U�ϗj	I{F*�]	o�p�-�߳��Թ?�"��b.9���u��3:4�4�ӭ]^����⎧*����ρK�Y��J	;k�pӡ�1�ѯ��>X}./�`~	J\�©��Ғn�}�l��D@q'fNQ	]&R�^��E�1(q���L��@�\�W���s��=~e|��l���
Δ	Z�����ؾ �L�1�!�n��iA�_\��BP��v=�K?L)H�譃�=8ᖈ���!pyn�
�#Z��a�Lm~7�e'��s��!�4�D����J�?���z��>Cj��9��W�傁X�Q�4��g�XF��?r�$<s�kt+ʆ�P ^�~B;шp�Y�L��h3
��^�l^_ ��L��:�{�xx��/�!��~��1}�9�>��̱@��S��X��M�9w�$���Qf�BS� C�MY��qԍF`I�Aa��l�'q7���U����sb��Z�����r�VdW�O�)o���ې�������E}�f%HXe]�M�~�~.Ϲ�������{���6�G�J�cyX*�����;q�<�A�.���kvL�d���e��p���l��!�
�햞��U==����V�]������|�e%�1�5���2ք4�����
����QH�)&]�z0��t-1c��c�-D��0��J�G,ydyo>hZ��<{���d�'7��K%�=_M��Eׂ���ڷfp���!%OxO�G�Ja�J���G��i�Ͻ�>�M-�H��0��[h����]hg��Өټ6�yw4(oa�/�Kt�=d�#����:_9y��S���)c�BU�\&�!��gp���g��{���	��|�~��m��'�������F.���wh���Lg<T��378OT�1=�[��7^I~��(��[�=}���Nf`[z;ٺ�jR�0"�9��9i`0\>����7r=��XRZ����'2��+f�؎i��r�o&[�_��T���p6YKe4��Գ�_�>41�!�:���x����X6,��h����18نE�ֻ����(5�qӼw�`BZ}�<�ctI�I�����H�L����b���!����'e\n2��B~��9:���$5�?<��-#u V�1g���Y=��YH��?�*i4@�Y%-̜UW&:]���O&n�~n���xt��=����'��t�,�r��x�<�)h��Wk_i�4%�v�:멐�{�*Ej�h#2i�wbL2�r�lM�i�Ӵ
��'���W��B~?����8*��CI��w��|B���#re���!�b�&K1�{f�A ���*K��g�PiFT��ɸ��9"��\`)�4
f��nn�pM��t�c4�ʈ��j�b�͉�f	J�˞�[�c��P5'���UX;<^V��B���N�;�V����O;T�Y[Q|dD3�����G���}�^TYV�?!��*�y1Ǝ�bL�8z����٨�$�lf�Nv{�c'����H9�'$ʻ���Ϥ��0c�X?�|����y��?�ٴ�a
f3��Q�dݣ�����_�;�,�cb�h������Hg>N�ڹ~t����X���%|Y�[��������]�c�w��σ*7~�����P'��,'�Эs����(� ܫ8`U'S]��bC��k�1Y,Z��]��Ҙ3����-�H���Z�j������ �.`��e~qH&9��>g���̟�5��Q��|���K�S�ʇ�K�Z.l�[է�]_�.d�k"��2�e�8�4}���"��u `���DǞ�?.��Ӭ�=��Am�[p�BX�#w��&�mfҧ�m�z}
|������4�?�f�G�bQ}�t;`,]�U*+	I��)MQ�k�*���}��Oj�ͨ�x��}tp
r��ld���l*nO)�;��]����0xo���_ArqvGl���Bg̻�r����lh�^�l��7d5c������b�W��
6P#�S~P49���|f���YI��v���㢾C[�:�>���.�WEaL�͢d�h����.��˥�
#͡��L��z� ��	�J"�F8IC�+o�+2�~�MD���4�s>{f߱E�W�D��Jy�m�G4�U�*UgB�L�I�ϘN{��E�?.uz#���K><1���G/���ۑ���O��_�"��lW�n�B1��U�j��x6cnj�8�@ ��E���0��E4Tfu�s�����}pyvQ^�4�;\=�(�H�`�d�>��`��$���[ QjL-r[����Ϳt���}��Y��2�}-d�tд3W�ַ�q���(`��f0�.�u��n��@�3�޹X� �#�9�P��<�=P=]H%k7AV�l:Թ��q8�I�/�}B�/x���q���^�I	��ӗb?凉
RM(`L��&$��g-HY�F�1�����s;�L���]\�EfM�vX��!����ono��Q�ŉ���d�1�L��ob��Ҵ׷����T��/�F_U-�̄:��U?��iv�`�gO!�����XVK�Ф�H��zCc�N{p�Mm��8@٤��x��"�אY��3=������g�\��!jٍ��q��FvmD���'h�(T���}g�/�ҢT�+�I�p��B|+��t�Բ:���J�Rr�H�<�럋��x=����������<���޽(_E����1�0��S:d���Cx ?�3J�EV�NE��!��`�<:�UO�,��¡�h��6���s�+x
 ����D�%tPM�"T	��`�����εZ�qT�o�:03�ǯ��Ԁ��*������=�ki���g�Х ��`�wj�}s�n��R`�"P��R����'���M����ji��(��lB��=W]��G��!����r�<2`��c1���FebT��?�ͣ��v��.Z_E-Ν>ے&� Jac�s�s԰Ē�&�w� �R|�W>h���Wy��/���
KV]��.�Kt�x�I�`q�ۥ�C=K
�{*��%�$�wrN�S(����Y���Q 30��a�;�[�/�-HP��Iaj���9�CUM�}v��/�q���:@�\1�k�L���悏P��`��;%^jHs�M�¤�p�39�9�F�������̞2N���z�t���0��ch�Ԟ(��Yv��M잟�F�/�t甸��ً�2V���1"��> ������-��;K�3C5Ƒe컌f������e��(�?����ǧ7K��LhO�=�&tl�><4���3�W����C| b�:��_q�^m��`>`l�|�[������
T����d��n��c�����I�KR<��rmz�7c��AY���W|�A6��o<�9���	����rI���*�Ȧ�Γ��@����#=/���s_#̢�2=^�Ť?h�Q���d�qo�2���t.�2-�9#}�#��ż�}�l�h�-���:�&8kq�BT�(�X�=&z���{�-�5��g-��o4�k`^J��U�>�㷻iZ�����-�i��ꏶ�	�ì`L����?VZ���n�,y6&u�H�7���'[;�5rp~�3k�](��v����k��h_�<��r2J_$ot�� A�_��L�oMGB ��Cȿg#�����Gt�g������w�/)Ȕ��L�J�ӓ�ί^#��0M���H��}��[�]s����@u�c=+߃����̼�m���хSQ�|L�zHP����u���ۃo����6�n6���ɝX��_�OT������o���Hf���׮�����J@����W�ФP`�0�O��v�W$�  ����.�b���=���K�.d��tu/��܄#�����f<�1	?,����S F�z�?o���O�=�~U`y�Yn~q�@��|+��!��w�+�,d�T�24D�2�,�������	vSr�����޾��y�t���yx�P2�$x�߫�`�Ƈd�����cv���m��,��0`��Q�۝��� !'���Ψ�J5����F����m��g�UˊU/t	�.[�����{w$���V����(@J2����6ǜ�Ȇ
7^P�6Kp���xY{�&�,]�Ԋ�� ��$����gp��۝S�e�
[�F�E��V��3�[��I`l�t�w�6��R;�Qϰ):a����'���U��[d��]�M��!)28��7��<�DX�}T�P��m���-�ϟ}^*  ��]"�� JGK �c}}cO?f����b�t��#
�5!*�	M�Ə~�&���@-T����M�]}�a�F�9�H��:!��=[d� ��g$�b�-�ڳ���N��:�ʟX7��%�V�i�O���v~?CH�9Y�$8 +�MhI����OV>�D` #�l-!�^�D�h��s-~xpȍ�J�P��r�W��2l�m�Ae���*��b!���7�����&�s����(Qo( XR$�5Y�O��w���L���P��
�]J�����E�xE�^�B��^�_]T0�e��6-,V� 5j�g��OSD[E�*��(U+8�|0��A}��I�1j�q%*O�?���H���єs��Vu䵶���g��_�8�Q
e������Q �"���A663���!!e
��g��M4|��泄�Z�g{x?��-��~���Fo���%�+5Po��(y���Ǡٛ|�j3�<ʮ��zH3A��$x�u1���U<O�x_�=A�\0�;��Gj�����.�0i	�2)3�z^�0�"���ؘ7Jm>�+�* ���{`�Z�_�+eFD��`���r&�f��a������B��S�f�q���ɟ�ͅx��}R�`?�M��iK���X�C���`�X`͊���:��7:O@�Վ�,��*����R$�2��!Zn�0R��r5&	w<��"w�!�z[3HB�y�Vb�������2sb�E�5���0�}����Z#���O�"��{���9m^'�3�6lH�5A�~|��ܟ����s��y=J[��1�?�KY� �\A�����F��Q���r���t�]V~46C�1�)��뷢Wɝ�1�l8���I<��o���V�EB=���e&�j��#D�c�&c��% ��@�����P�"��Q��Ȼh2���,�SX]���hh E���U!���b���(�-22}�dN�c�)��YN�
Ÿ�m�xkyG��-�0�;#�~
N��@�݌�S�������u%@���B�x]��zI߈�k�cv+mm�����!ކ��lقr�݋Ru�-l�W�M��1$���R�(�b);���nc�ܟ�3������3�-o�H�Tk+@-p�;�^�Q��$A'��b,o��k`�u��:72�*O8m����h�V`<I3��K4$�����ƒW��&%wC{T)~J,w���`ҁ�]~���TYѪΌߑ�;���4����]hD�.�Dw+~핫��]xeUi:��t�DR�b D��ؔ�:�v�V�J�/`@".���j�&�<���kT��i0��;|�S�R^B_F��3ҟ�M���]<�U�Z�k�[ESWJ����W���I�WnK�0���a���w�cRN�]��]����3gE�~�똴9�P0����*��0���u]�� Yϣ��4{�">�MQ�B��z�b^�,8q��*%iN��C�ZT[������S$=����d�uI�ޞ��xV������km��	�ۢ\�UDT"���H�o�80��T��P+WVj83�Ӳ�����=�P��FV�~t�p�K4Iy�޴KC6T���"id�^Wf���/�Eݗ[Go:-pr��;�Dz��n��HN�g$1��\L��!lp �v	+f��Y��O<6��To�Vߎ׭Iڷ˒��{A�cN��0��Y�I��?#^l�ߡ��+g[�>�)R��r�b��3S�R� �W{.2O����il�������6����;�s<���i���ڵ�vv�/�]��?8�류�k�V"���� �������fȏQb�� 3�`ǻ��KI�Մҁ<�i��"��5|#��q�Z<Ql�J�>6��Y����1������0��w�'��p��%qG0�N�Y�G��Z���Ƚ{�Ә�d��I�GD�z_�x�h������ޏ� i��9P)��L}�u��Z���um��w�:`OQ`�rL��S��h��eb�I�4��-�l}�ٲr�ș\����c�h�;���I����}��W�/��|D,0Ug�lsK��'OIL�(ތO�7U2��F�;�EӍ������8N�V�e�GZl7ԯ�/p:<���ULcF{��  O7��`��3�On���| =�m���V�������iA+���"���q��������g�ctO���-1+~�#��y�`3Wa<��|Y��=h�4�� (2��0��j�Fq���4#xK��V������NS��wldw���,�����  Hx��^��$R2�!����ҧ	!���A�i	*q]HqJ`a<v�`_?C��i.Vi1_"Cݲ�<ƈ=	9cP�s/	�,�1��#3��Z���,H���"�H�˙Q7Sk�H�]�p��i$�$��KZ���vku������X�ޛɛ�̷�(f��}��F(k���ç��^&�����<�6WKWP��|���`�Z����G�Zp�Ι��):t������b���Ɉ'�� ;;j���/��q�f\��%,��F�*u��0+D���t�g�ɥX�Z^� +�B5��<aY��#��.��������\�&�*�K�&]Iϐ6l���n��v��b٧ƌ�k��i��^�����5:`�t$Db����ɖ��Vj��+�j=,ܰ\�2*X���Z�X��#G�O����TI��Mbqb�������)h��J]�W�eYC	FPjqOx��!'@�Ӆ���x ��-N)_�Vw=6Yu�q8.Y�WW�����\̤W�Rw�� �>�=dXqY/#;_Z�O2����K k��!\6�7� �(F�P�K��r�ToZR1�HL�i ��}c���h�ߠ=8) ����6nb��O%���Rs|E�1�m�.�O�7Pj/����U&��!ϫ� �O6��Oh�2�z۰��(=�, @n�q!�~e!v�:e� ikc��FX ���#Y�����Yx ��׵y�m��T5#�6�$�^@��IѴ[�较�m�t��]��~���l	��
UW1E����?4�7S+��y��A;ߡ�x�6me,e�I��OE���#��=��7����Et+~`�I���l�و���?�L
छQ���
�%l�M�"f����T�v(i�~W��c�;2�f��3�A�mR��0�F��4�J�$o�\u_5���' �>^�2�~�?px�?��P7t���$?���u�rv��y.a��}��n���>#��(�E�n_��?Ə�k�܈4�"�ܝV��**�Ă�ԡ'�^�D�d0rS�[�gR
��H���[� IM�<`�)|��N�>��)(Y�-�Jǚ'ͼͅ5�T��`�]��45C�硅�f��/�=�iN�{mU�h�n����ɒc�?�Vw�DQ��q��ٯ`�\��xҍ���`���N��	�R��ͳ��$Щ�o��E��)�Jonu F�;��2.�����I(i�`�WΜ<�_�j��ⅉ�ҏҐ�g>�"Z���a�=�I$�<w�z�@�m���_�¬҄���|�`a�W����GQD( �]i/y��f��]���K��'��G�!+��%����M�k�
�ʟn��x�Z��Q�JdLa�@�N�˧�����o#��i�G%sLH��q���q)ghx��d物��M���nߗ����Η��z(�;�q���e�	g4c�Ӏ�b��+��YM��d����m=غ)��q�3잸ϗ\����j��Yr�nR�;�T��U��0�sW�&�p��R��"P�g�!1�'ye���Z������n-d3A�`��yd�I�&|�Xע+ڢכ��J������-� {5-ZDNOzy੟D�/G�a�r����v@�ͮr�M����W�pAӴ��;P��$K����A$^��7gGɸȈ��w�"��2"���� �}�u��{��I�5"et'�3�Ț����Ă�n�,/�5�K�A+����s���z���﷜�$�4�z�ɛ�FZv�+���tEr�H�(�F�Ys ��
�*YNB�F�?�m�C�޷q�7*m�՚�5�8e�&iŹ�G}I��<�������,J-6 5Z��1A�X���8x��,�߯H��^���I���,/9�����aac�)�����UY6e���n6B����kc��2m���I	��;���6�,:�>�2
EԁU�<^���&������5��Q��Bz�W�*���d3:���{�;���IJ�����RG�7�X��w�45FH�ϵ�r�n*���&������ u�	�=ӵ��z�y���G��\qX��n����ώr����6�g.&I��jl�]��j�|y���P=H�X�:����;��XL�u�~cP�-3`���[m��ͥ�>�4Ad��M�J���tIسqR���g19`��j�cW3/���X����B��|ߜH\��ZX�vFm�f�5&�Ʒ0|6�z6�r�ϸ�U�Ɵi�'�	2H�w�s�Ŏ�CQ�W��l��SoTl��{�"4(��{�	mC��|J�g/�ϔ6'�2!CtI�Юp�r.QC�/�����E�;[1�ᡤ�U�:<�����D.o�)j�"��)ɧ��NW��e�Sb��e��	�Vב���A�_�U"�=@)P�xC_"ITd����,XM�)��J��Z����Q��R���F1m�	Ab#\O�7O���*�xV���DCRy��^���ou�ǁ����K��%�[���Nz��<5Bk*8O�'��	�V ��q�={���j0yWO�r��~
�采w&+����V��D��	kf�o+a�C�R��5���Ä�>*���k�{ j� ]�	��2a�^���Rt��A)zO���މ�:����3L�|��Y�T7y���� ҈M�fg�q2d�'���1��UJ!��;���6Mk�j��Ք¼og����Yo�e�\��#ǣ��.��2�G�n#I�m��ki�%I.�B��l�z+��4l�#���g��U`ڱ�|�l�G�JX�R��;�x��cڏ�btZ��}'�$O�@���t���F�����a�@+��>���?���� �))�L��{*�+���Z4��bg`�b
��
E%ʍK��&9C���_�Ԕ��va(�\P��M�L˺������@25�uA�{⦘�C�s�~�:�O)����c���� �2���nj�q
���
w-�mz_�8�5=�vFJ�0�He�L�T�Q��f������&@w���;���V�X��M�.��H�$5�����:��W��fT��Z1Xթj+��Kؐ+ީ�q}�P0F�̙�&�?���j�0JC*WC��Ð��h\A��r'W������k��nFN癰�45�õ91N���y�Tk�xMu�D���oz�����y<5�ὕ����"}��8Ù2�<�͸��G`��mt=C�RZX�>�M�9�$�
�p�v�h+�}ˎu�	����v|�C�	��[�K�e��k/g�9�V����.�������遅$~�Ъ�|	 ��b�%&٩�ku낱�u[}}�v�8��V�WYV�l,@��Sl��u��nYc���i5��� c ��~[ԧ��:�g��Sw㉠9���(�/;Dc�GR�9�����WԾ���H���P٤���[�� �~rd�u:9 N^�ED��q˘v�]Y�c��k/�~\
��Xn�!+n2Y	/�4���x�d���E��
JF�\Q|Nq�����Ng�<��$;� �=�K�{�Du��0�Jx��?=��b���>�+:FK�M=����Yb~*̰?�j��"E^T �aa����x�Z����<�p�iԕ<�5݉���צ)�ڻ����Is�d̎�^3�+�V�Ho��RZ�v0>ۘr�@�ٓZ������"��ʚf_�M���O��7[6�R����:�F��~��O���,$�ľv�۪�6�(ǂ:/���}��2���ҫ���5C�>�Ԫ4�h%5`�8QY��eD�"��]�%��D�\k���b��pw.!�e�b咟���Ҫ��x��U]��<G�Ί7�,=�j���UΐdapL�/��Y��dc��֗U��!��D�j�#(�������E���́#̡�zA�G|V_[�Y�'mċP�x��\H+5�	����״�ы����z�Pp�z�B��QTB����e��WW`��S�!g�@*��bm=A=�Frf�����6͇x�5�<��r��f;`���3�������,���e�k>P�tDL�gܩ6�sm�ӿ��IU�wi�TN�i�-�A&~D�Vu_,�Q��~�	����8�l��E�R��� �}\���\YJm�5��V%���h��� F��c���#��l��0M����!����}Z���X_�՚��=�Զ�ᯉ�� m�}���z��jK>n �4��=�q_���z�@�K ��C0ny���e>�K���dz�M���n�ǟh�y�� F�0��	�uXa�:.F�zkbK�Ÿ����X�",]p.K��:����i�"���&] ��[UWE��o���%�v�R��_����8�q���t�њ'��;�Ȝ9�Ow[�������t ���&�o����y�w`�8�j4�4�s��
��I;�)X���HZ��u�C�쳛�L��Dp��ө��Eޒ�m��צF�<n�(��Ϝ���g826���,kh�ͫS��3��ڜ[n��Hp���O�hG�%3�ڲ� �������w�*�R{�$i<�t]Qي]%a���?�|���� �F1��hqn���K�)�с0T���=�"F��qC��풃gi�3�a�3���iĻ�BOXl��WY`���nCr�jw��x��G)��ׅ��K�MfP*NVT1qN���i����_��֒.��0�[Gt���:�[��Uw+o��^S�%YIgP��k���w,�N7g=�~�u�z�mj1D��q4���i;M�o`Rj�&U*���*Y����H �@�i��מ4��]k� � ��w�KRth"�P:��a1+��}a�`�E��R2
��B�~���m;��d���q^3q␢��o�lW ,%��Nb���.kzڃ_љq��:.O�b<R�d!�i�Z�ˠZn�<݊�˅J���X�l�Q���E��d�QMI�vyh���Q�c�[�\*�N�Q��N��� Yk�w4B�����"}o<y�yvA�!�X��q�̓ m�1�	��l�;��0�����f�aS�Ԅ�>yҺ�=����3����O8��o@���CK�����@��º8�1��0�P8��/��[��� kR+�Fr�/"��� ����P�&U���Z���*�G�.q�����,Y1�Z�6Kج%K&��!�H�������k��B��M�g ^㎎Ɇ¶���������fE]D�&�vR>?Gu vO��ݐ/mmZ���_�:I��������Xk�O!'��DH��h'��!Ӟ�r_�7��)��<Dp�Xy��� !7݉�@N5-���f
���bb���0�A�r�0`a������T䴽\"��mP�9�P�~ �ٰL����[����B��ȣ�C�&f%b��Ģ�1#����K�u>Ӽ��ћ�{v���R;}�>�ng_sQ���+i�?�h:^�����er���5q>���cؗg�5$NNN��}��]���^�NnȒ��i@��(\�fZy���
�|'PV,u�ۃ�btЉ�i�m���m�y�Ĩ�:��^�.���8����M5F?��!�zP�l�h��Z��e���\����^U��#�;)�lb�Ze�LO9�.EZ������_��{�{�<��4-�.^)�l:��v��Lb0G>�m5���`��q���r�!8^ϒ�^��ZQ�C$X�6���QV1g�gl�(]�X��8���?��m�+%-,H�	[���%���p�ً�|�ӗ����U��@M��;�冒9�Cg��{:���d��l��jA�7<��4o��G�O���kr҄v�����0��ث��!)A[��>ˇ�\��gf���'%�����BT�X 3�����e���ՠ�!�9Q�n�-��01�'����%�u_���"w�<udѦ�����v�ʩ�]<)l��5L5,��X(p��-�̍�B�3��醏(��6���7DMW혗�=��H�v����C �O�E�LIW�$���Vpee4��;��Կb�X4�6�Ό�Tc���8������z�=�"6�׋�>V�޽�R��v(�����o�MP��B�[���C��$W��nĊ�	Z� �e�1+ϳz:.�s%��-# ��_���b��D+���2�����%���J�>�m�X���'�be���|!�T�Z(ySK���}���ZϮ<VJ�ϧuC�o��-�i��
=��/���Aw��:����������K�}ދ��rsC�Ѣ/|��p-(�+�F|u�\-��-�]Ȃ�1���-�	g|��A��P��.��� �z�͞�5\a
�'L/���B!�k.oo�1 l�Ր�2R�`�@">���t�|-D�S;���b�D\B��[D(1XK��Ā���`��^�-�	m�5gt�٬!䢦=��1=��-����ԁ75B��Eۣ��VA ;�&�����a�-#d$?��������V:h	6�\ݱqȰ�'Շ@�?t��awe(��x���v���^*�E�~ )>]hfU�Ӡ�\�bu��T��Ʒ}��!Ȼ]Kf=#�}�]㸂��$Ț�h�C6��<ܩ�q�b��f��9txu� ?�F���Ȫ|�����p&(	�Y�w�8��{v6�;ΌY�jO�x��+��K	��Uם2�Ӥ?�/��h���/!�nP�VEg�h�w��V ���%�o���A�ـ@����\E��CoZ&���&�L�&
����=R�+�k�寁r�"TW>)g��Gq*]�q��y�bA�f�����J�� P�G}�ҷ�鿩�-��y�葓�c��S��>Ky*R�f'ҎK�Z���2��h����K�"����{KL9���Y���c�]0�+��T��%<�R��9�f�u�������hRU�� �l|�%A��e�z���,���A��	��,"H�CB�����J���x��Ѡ��uA���AI�n���"�W����� ��c�/q�4b�q8�]n񬑖�3l�Ԉ�U5W��,�y����Wx��jK�lF����q'[��⸞`e0�Q��D`%^)����9���H�Q���ρli/i����78_M�|A��>&��	��Y�(S@��2����r��J��&�=7}��[�d�B����1���ZΫ6ڜ�~S}�^����?�aq���<���GIB�2�^l�bɳ	�$<�~���� �Z��R2���*T��6x�6y<'�AVa�ܾ2/MG��}×���P/�S�}�Ml���#��g2�����^���Z]\�}��>XHi0����X��Ѽf���n�U"C\�;�̦��oW��J�Iv���F��l��V&���=��W�R}a~=�ki]c��ly ���X�#I���'�,�e�>!���ePS�4,�o�iɽ���� ͖�vϳe_�S��L�HA�F��dzb85[{s�����D�7����CE�.�R�gc�4.WWۈe���1q�$7W�`�����.up�6U�:��b�\=gz�4 "#'=C`R'�9��$�Z����޽ȁCpei��}����t:ïM���iąy���^C�٬�ys�mqg6�FG:�+��i�����B8���]�O(�̧���F٣T�%��$�v��S�D�<��-6VϬi4�`*�i�����V���³t3����w�R]v�aq���< `�|��m�%ǜ�B@�w`�1ˮE�BJ��M��\�\�J�}��:�����~�%���/��Iԑiۤ�ⱛ�j�g_78�7�]A������e��{2��8������u���fp��S�fN,�3!C}���>����V����)�^vS>��ɷvoi�g	@�T���-��zI�j>���r�df�J '(�`�M����a-Ę]��w��)�XGl��ܥg�b
���-0�N�OV����{�^֥�欋T����	l�>�qZ���Cm��Ը�Q��o�)_�4'*���V���4����Iϑ�1�����)"��`^���T֊�ܰS�\�����w��'�~ŷft�h�<J �gO	y�M�a堕)�G�='�gߺZ�&$�v�J��_���%!]�`I%�,�8��e>�p�㐉?�v��(�L
#�������t�?�+v��a���[P7t�+�s%-( P�č6�
�vA����'���`\�7���U�#vz�,���zl�[Ѩ ,���67����e*�ӷ^LP�M�峍��{�.��� �p�7n�tp�hbjԇcjvº�#u@�3���WWkk^�3.$;ٙ�4[BQ�I���w���m=��e8�-T���f4'ի�?�����_	6pP�ν�Lt�����L�+#�"��h8LHr"��N<2�m`zM��r�{#��_h ��� �Ϣ��$��6�z2���C�>�	q�Kt;r��vZ�Qt��K�7)���z�&��W�e�N_�����dX��;���/��;�Ƶ�Ls�,kg��vM�,);�a�Fe[�d�R!���&��Aܜ��n8�tS��8`���`k҅'�b$�;�0ڑ�B78w���Q�qK�<rM��W��v���6���!L�9��-���x8����H�#x]�b�(s���|:�8,lw�ʿ%�Q�. ���L*�S�*!�5�Z���!�G�>M"���i�
)2u���R[�yo�A -#RRbz� �����U�'}_���Dh0�X�`���x�Rcݫ5I7�ǵ���̧y�#i� zLiv�.���K����_�L�vg'�Ȱ�L�UPF8�wבf�]v0��	�6�
(�����(���LX�w�Zcf�g�|�cA�c\� ֱ�De+F�ǒ8��0��I�Q�H�sS��$x��d�@�����%��E�R
쑥��񘤗{�<�p������B��S�;|�Ī���3N-��4���a?��� N� ��~]Йs��a%�����_��-m�/���v��;B�sO#�p�Աއ�.%�~��4a=��uSVS�����fH��'&Z:l�����E@�:�I�R�������F���p�(���/u��z@���5��@|�էp+���̽Ÿ�%�r�󂂪�d��h����ӧH{�%�6FWr�k�T,o"�����I�2�ݭ�ܐy�e����_{�5S�v�L-��\![V�H�3Kb.-����0[�O�2[�c'�d�|�'<�ٕ�j.�b=t;��Y~G�o̳��%~�������PF�?�2���Nn!o
v����FޞR�ś��v����Њu�3���)b�o4�����YKi���q���̬neK&ޛ�|�r�<.�$�Ug0���]�s���w�fxǪ{�P�<^q��?eonW��>,��v*�f��ߌ8k8�A��T9�����k{���O-a�?�>@�c�g�T��p�b;X�h=-�
קȾuK�1�A)�Vv�I��M��-g2/KL���t�0�ɓ>�*�52nK� ����J�r���9,�B��*�Yn�� ���o"��3{��O�2��̌-��i`U����׷c%�L"+μGM�;UG���O��N*�?\���2W���ƁW%��+�<Gqz>�������P����u�>���i��>�.�ѪN�,"MM�V?�{���{�����6��2E<��|�!!�����q!�{�I�_�>_?N���}��Q�����)�H]�o�6*0�u�B�B;�$Z��ݮQbdQ�}�[�v`�i�/+���'M4_+IJ:*�\�KwLB�M*��3clҹ���ÞЫZ���*�^��1�7:����0�b`�����`Y�xf���@G,���x�I��E�q��TqV��a4�.�~�.�5�S�c���@�,��˧�-qk6�ؔ��t�e��W-��_�9	�P��x��˸��`x�ca��s�_�~{ڂ+��l�<�0UJN�v=���
T�)�T�0����mS0�~M��Uk� ߟr���
E4�eOߞ`�³�ᜭ�'��7>�0�r��9T�U�3��C����w�Dy���,��'���C$���72kxT6����nDT��ag��<ȝs?���F���{$:<P�%P6�^�1H7�rЁ�xZq��A3Y���5�$�
q�_�R�Е�k}$5�)�,�9wE����Q2�!_�����o��9g��'���`C�P�8��i�M�v*�6@��&�z�69y�JWv�bL_��n��˧=��H�}"��U����e���1�]ɓ��e`�o�Q�]RTZ��Hm���z-��@:�#7�C�[=j爫�w�Cxճ�'�ei�|Z�KqiI6������l�f���y��[hن+��#�y�% �ٝ�`�pU�
jPY0�/�̈�E�W��|�:�=_ܘ�5������פ��r\����5���xϯ5�O��ۘ�wٹ3��C*����嵦��KU�Op��)u�<dt��W4���$a�z���J��y�[��0��S�� Z��< r�M�����(;߭Iʗ H�!ھ����j�عY�.��](o3!u��ZP��<�7��dd������3寇.�᫔��1e�>�����K�7*�o�iP�6�\�Rq���~/F�}��h*��M }n���x
��e`�3�\�B��KC���{�xw���`vϲ�p�<��|�I��흚�ky���1=�e�~1��'�V�)z�ѧ0pk�TS������ụ��� ,��Z���BZ�l?��L��7ғ�&^��785;7�vlC�� Rmb�ݷ7�oE��P'=K"�f��1������R�U�i���S�$���۔E٤6:YT��R���$�)�B�6S��T��JC�Er%N2'�uO�f=��0�<r4�|=f��̹�%�u�y�Fǝ���2�@���M�1b5	Q&��\d���Zt@�F�.�Tκ����Ģc�l�&~�pmI%����&��]1��i�$�$���#U2I�������h��D��s�.V�	f8!�]R��]�E�-my������*>f�ʪ����l8'�f���
�3~��:� pIŇB.�HnN�8��q$�$�8Q���t�QW!z)~X'\g�r��եSAʟ;���嵕w"j�j/6�4K��s���NG3az(�,�Q���3�yRF�m�F�naw]�ł�_���b���B�� ��y�������>���f�D�X8�z�$Ձ�����ᙡ�	�hU9Ʈ|s���j�HC�T���OWY�1 xmuƺ-���S����_��o�zW�R���V{�J�����؜�����q*.��1�XhUW]q%'�h���}��v'c7�P;w�<5)�����b��=�&��4��^����@n�𰗛;s�Az�
�"
��`=z[���uZ���%!�#�������;f2c�E۹.c�l���у!K�\�
��)��V�b6w툟����^x��i�T�~��wH����d����1\!tm�iػ`{s	�~��N���^�dٰ}Hkd¢U4�G��[�R3޵yL*꿓�ض&	��7h�Ex�\�2���{;��kZk�"��H5ST'�}�� =�o���*��n#��+(��"z�y��@�{�~r��n�V3�k�.�q���_yc���;zW<G��[�.�&oJ�o��P-���������D1��PE�o"``�+�ɤ�]FkoZ���O �c*Cb����5ӓ�ޕS��oJ_��۬�a����j�~J_n�f� ��J���Z����� �ΊJ���o�56{�6V��9���7
�uJ�/X��TX׳���tB@�w4��I �~�(|�R����1_��})��쮈g�6p6�����{�>�r�O�M�R	D�������k�Z��bt����{� %� ����UL,!���-̖߃U��)��o'9�nhS�>�J�S4��h^�wy-��o�jËPG�* I@_�N�{P�E�W`��p���}�Ƒza�����~�=�T�~2:���,�W�\��a]���=f-z��(�Q/҂w�TZ��c��O�(I�saC��F'��1���pɮ � V���d�R�A\��5�:�LV�������Yt$�e"@�7�ӈ$�L���<�6Cy@��(���A_��gh����|L�?J>�]���fg)_e�q�����Ϳ�{�䏑�9E���>�RuW���ˑ�3����ۯ�Xuӿi4_�s���򓚁3�ⰰ�-��JBq�mr�I��!�3��|�">&��)
9%�4g����k4�2s�	�:���'�t�MĘ��3bT������3�G���/��u���ڿ�ul@��PX�J���YD�;b�}���߾�|�0���=���ڛL��\�	+��%��~��/��إe/K�V�|���+�z+�%��A4�T�@�����-�/HW�v��KT�)�������"���;��/(\؍�s*ׄ�!���K�wW��¶h��x2��'UL)6wP���)���x{�^R�5Դ\N%h!Z
�5	y ��G+�i�A��	��L�>�7j4y�_h��ַ�WA��֌y#�t���1�����S�Fe6���k����G�תC���ڧT�p��W_=H�����[�~��)�2GR�}��pw�5[SMҐ���˞�Qz�{�ߥ.�E�$PkB�g��4JDۦS}��R�� 4K1�w�r+�"�z��¾6(�z>�ڌgʦ�~�nK�;�8�t��b�[w����ϨfZ��L:��bi�$hU��	{҆?���L�i��x��3NP����i4�,�>���)i�#���k2kiF2Ƈ�NcMp���΀8����-�\�I$�q����-x?���a�����Yhz��mhr^�=MԦ�u'���'���^o"ɑ�;�DBg�*ا�Z4pSx��pv�		G�FkA��%�z�~~+`Bmd`3�.b�Nb�t�^ؾ�����1���f�vv�B�2��5P/�ߍbl+%�k��9Fr�)},sx��@3"�)���ѩۣ7�> 5��y��xLMpe���RD�$X�U�Q�7��u��~�H�����QLwnb�
-��B�莺��eS�{N�?���hL;>*'�� ��1#�Բ��{|@�(R���(~�<s�Pn\*nN�-�դ���^�M���Ҭ�Y4+50a�BAfbxL?��pA������ɖ��l�J�t!=�4�N�x���q�-MK���V�P��������P8�DJ@��_o�;�[ḩ�V3j����`4
<$�_��zM��30�J��@}C�#���6�\���9��*�����p�hsm � ��.����ۋ(��|=�t�qŗÉ����7J��N��Γ�]�l����W=r�I��zpR��������cc@deC3[s��~c9�k�W��� �*�6�B#>!�����2S[�r�=��/�tw��J~�­Z��������~�7�*ݡ:X_��L�����r���jgpV@L��l3�׿��ٚJ�}�����c����3J�	p��b���%�8�ة!aA��w�<�Y�29��#|�[
5�O�l��u��"�sєw9�A%5��\@�O��i3�.���m(��S���yIz]�g̰lQ;WE���i�gE��ћ�0�*��-�`4Q�:𫲹��b;�h�y��D�ˊ)����#�M������{o�����{��t�ӥ��hY��zzx`��ɢ0Uk�PN�I$�G�C,�H:���6ZG�"�vq��Zߘ�,��k�C�T�H:i��_����▿�z1��1�ՙ�V��Л�|��h(U�n�CޑؓxdA�Z�&}���Rd��ItԦ��m��rq�Y��Ʒ<F"�Q��P����wU�G�$��Za�$1��Z�%���sbX�'ɂ�� A�*�jb�ڴ\��K�k�	=:�,b�C��}��#��iV�q^ �&4��R[�8�!< �6'����TRY6:��_*��W?X�[�*���Ng�i�KI��_8ʻ@�M��9������*�	FX����|�F ��{0t��-2�+�M�^�S�-l4����^��S7��4�L;�{0Φ��-���eGn�~��ԌD��@��;j@�S8k����X\�q�ۤ�8܈�T�ێ"� ?j���Q�4��B�\���|q�)!��B�48��P0���I�s�hzrWK6�(��}
&.R��j��椗[�~w�H���G�^a�&
o��$f�[\��B��2���s��K��8��|�3jE j<��R�+��y3�u)ma�f�;��x��o���0��)��z�ࠒTD�)ԛe�-��^�[~�L5� Vp��Jʑ�0+�Z,>�K��Xt#L
2���.l�-lF��J��)%�,W���_(����МhK 0|1��"!�Ǌ=R��c�ډ�^r��A[�+,�Y���+l]rنlHʐ��)�� N1���ӫR8�gd�:���R��gs�$1V�� ^��M��cra�#�G����!���NXr�83�Gʠ��$B�a�h�������>����~�7C6��xkh�ni��co��ۨcʪ���:�l���F<cP[F����}���g{�M��b=���� U�,ˣ�*�\O:�ݛ�s�Jޯ'�]m}�b:�q�/�YŪ�Ĩ^#w��dF�q�wOὄ!ypK��ZE��d�zc�ޏr=�]��p5F:���ƒ��s4R�
�w��������� �����L�e
5�$�1,n�w��ݺ##�F��PD9�3�i����Rf�$8aoc���Gp�vb_`�Y�Ü�Z�:�HjK��w����z��(��U�;H���r�ـ� �=%H��گ�ֻ!�}�y������֝:�B�K�S��
��!��Zx�C]p��w<��8X�����YNK�LA|S�J�'؏U'L����е�^;!>��㖛ٳ�Ȟ������F���Y��2��!���P��U�������?�	"�����S:�(R���v�nD!�6�)�j׋��G�xj O�k�pz
}(�rQ�@��ϟ�p�9N<��q�F����$�C��	��������p�5��K� ���@�FZ�1)��+̠���ւuaFL�J��!\�wz�btM��f����D���aDw�Zs�d܇�ʪ�C��F���h�&�Z�R���<hM��2䗹4@M���&��<���>(q^{_�)v�t� ���vrY�U�#�`)���L���:��6h��h&�劀Q�p%�~l��ԅ@�;u7��W�'J{���P% ��G�{��H�)����g���x__��$��Wp�#�� T�c��(Y\�R��M��(*pf���������+�S1�ӹ��j�Ol���a2J��
����͸� �	�z�x�=
�Fҋ����)��=�j�p��T��xC�q�8y#T��ys�hq��5��pH��OK>�'2�t\��2{Q��%�L�����V�����JZ��}Fܞo��'�yR@逝�p�뉠����U� :�a��So�}�G��i�w5�F1�A���В�o��!Z%�8�'>n���L���FV �9G���ʉ��m�58;���;���
��t.�PN�tXX[&H�PZr��μ�Ƽ���I���*��d/�V���g@�0�_�Q�C$"}�ړ3�Աed�QW�����ѣ%>�9��>�!����~ò��z_�����r�Τ�lOד�#Bv�U�Ʉ�w��V�uu��4'�|�<��ދ��9��a��H�{�l�Bؿp�k\�~y+Q��6�nMA��get��t�>����:���L����gn�"S��Uۙ�YH�:F��N��>�B���Yi�l<A����?b��1���5��/�MU���k�<bT2Zl&R!pa����5µ�ܛ�M���[^Z��${)��P�݆�\r��\�[&�d5:�R��}�K�4��% �K���[��|�%`+*Z��i���/2w��}Pd����3#D��؆����혢�>��fP�7�x�;\5h�{�i�޽�~lV�vK��n���F��(��7֬�B������'y�QoF!�?{�2q���뉳�V�4d'"{�Y�'��W�K	P�'2���8]H��x�8'�'&�1�A�?��XǇ�m�����EW����^jk�1�2t�0���ӗ9��|�%~��+
�땀���_���ܬ� 6��3��N7�Ɩ�����ǲU�m��Y$�-���z��Mp��v�i`��vڹn�ۚ�Ax�}�LD�.0�~q�?�T�GV�5�zT6n�H������]5N�����|}`�0����r~�7�[��C�n�e�.6$wy�o	���n��/n��L�KVcAr*V�4uy�+���`��d&����9 ��@M�^�������z�6��,ҿ�[X��ǃi/dT�3 �$H��W�%>�Oàiq��l]=��E�&����z3 �����4�.�]�?WF�Ų_��u
���)�BYJR� �!����(�/H0Ud��ny�q���%�L1曩E��3�2��g>1��\�XEZ0UA�r#^K��Y��淐��򛙆���� <�=��\+���u�ф���O����㰄Ϩx �X 	��m��ҵfqz��m�0�����Ѓ'V�I&�y����G�|�A����@���t�)05�P���
5д��~/<��]>��ؑ�;�o��9d��%ՙe����.���<DL,F�#u���Rd����qR�=O�x	69�mǋ.�� 埊�$V�/RnMl�����A��xꉍ-�,�@Yw)^c�1��������`0n3�A�čkx�c�����j�
OHe�Σ*K\-���o"���o����"r>w�2z�Z�΁c��������@�D�p?�%�;�I���n~$���,��x��&���|�DE��ֺKF��A�P��
�A<�#��׉$����?�&�GN��QvR���M_��[9,�/��s��2;F�l�����Fޑ�а��M������l�`���.N��nϮsk�w�IB���/l`������V�T�z�;�y%��4"��jA_�n̙���4�+R5���Ic]��Px�u��j�'/+w��c6���T��Eg��g(!�/�0[�6iE�2�Ӗ�rb@BH@4F��fYz�ڐ��@F7��݌^꡹i<��N��v���b}��:u%*�i�2-��|���x���a�z�{�E-��m4�{H�nq������^��S�ecP���|mQ�p��zG���	c]hW`C̚�M"�@w�Rs"b�_��S�m=�cH�1��Y��0��+N ���NR��⸻��Y^���%��v����|��u�2�ya|�]	��ǿI��w��)mss[S�>S�绰�T�������$i�Bp��V9ٳ%-�X�"pD�Q��Ǐ�qvܢ��e��1�zm+ "���jOǜ2�C������Ӿ�X���-'6=����S.P�]��;���T�O�\�o��AM�/#K����TN9�鍇�\���t�I����o�0�)d���F4���9�x��}ą�B+����0���x`��v��q"�"��tY� �����9�J�K�!4���a���Zw��3RUD� #��馔e�<�&I��[�G�ɗ��a��tP��LD�-eO�vP��|rN�6YL/�/�ydU��d6S�:�a)HV1������y⃲�_�>º-O�N/.������_��Xc�@
K%,lX߾��������<V�V1{�Jc�9��e�	#w���?��&��A���ޮ5ܙk�Q�h_��{>��Z�s��z*�uAK~�����a�
��瓼�q���b��5o&]�.���"�]�
��s&�|�wZ�78���H��i�Q�I��ω�au��W{�hXo��-GѼ��6:{劥�I���	\�{�ݥi���u���'���{y�r�%�|���6g�?:t�f/�+A�Ѥ�L.�|�C�Db*?4���/�Q y=!&W:��*�H�φC����K�s#� �ʊb`�(����~�	��T!H��`e�R���jG�&�f�=���J^b|�����8:�j���!H��&E8P B9��8e�6Z���S�"BU�2j�.��owG�WY�F5��}�l�-_&Z�Ú�.�B�qvs��!0����c�1Y��\���`&��cuj�=��V�?W~uo(NɾP��&'�v4�0�ؓ`'w�rb��@
g~�r3����h{hA��qeI]&뵦���U�b��G�E�������<��G�ێ_�s��;erY�\ܗ��x���ںT�>>�gk�@���7�
���1k��od�ӽO�t�0�E��I�d^�W3���ulY�v�����3���om�F�
�b!�P)�y5��X�����V����;2&\j�Ν*9�X�����G�ґ�ʻ������d��S6��6I��`d#�g오��U�l��
�}�C���$i�k~" �@W�N����f�(�_�A��T��`wPGb������L.�IU��ﺈ��4Ñv��!�i~�{����rХ���fME{)��0�2�f8��#@�q>������x*VH9i�t/��L��g��,�H�/�$X��>��E�E��W��h_(|n����Ň;Tma-�(e;����ڵ*��^�m�˨>}�b��;J�u����i6��s90�;�jtXҐ���sr�4̂J�.�9��?��@zZ�Ő��y�{ɶ�er��T������_A�DZӹ�lҾ��%|Bi|^F��l�&����9Ya��5�mS��g��*��=�����"��ͭv@�z?�n�
�)�N.TLBV�V�8F�G�F�6�kppe������2�[���-�$��$ &�`�s\e��^-�nc�ߔ������sK��%��gZ�PE�=xs�)�.'	.Q1�#�D^�3����7p� ���b�����3�~7!.P���
m�E��ː����DJo{v��ؠ����<��|yn�U;�id�C$� �u�������w���` o�4����wcy\K����hV��$�Hw��O	m�B��s"��lT�c��=�55ɸd��IM�}�q�(�͙y���`
*���/	��m5�;m�U�)_I����mT-T� G151"��z�y��(��=�ypM�Μg��]��D��2�be��OBy��/n�DbL׍N�#U���5B9d�_}��z_�(���@�T�s�k[��>6w�`�|Ù���z���㾄�(&�,���������~O��v��>��_;Fh�r�\zq^�-��텯%�|�!�PXA|MPk�F�8/��iP�D�/'��	1��!�UR���?���70 KRy�b9�F`�=m^u��bJ ��o���56jU��-�C��b|9r��(O!g�U�0[(�ʤ�!�\��\_��@���d/�0�e��ł6;�X�,$��`�x�H�B�e���K�~�5����Z5(�w�!gg�Ȃ�J�/Y|��e���٫���Rᨇ�u���9���p?���B�����0w�9A�*w0C�C��L�$�,��pRsn��H��\��|-Q����� ��ԖVA�ޞ3��|��`�y"1e-شR�^K��z?�����􁖞�f���%�y��]; :����j�Dx,H��r���Ϙ#�7I:��6�rv3�`�lߴi�����o�J��㶭�Ϳ��ɟ�	*<'mO�9v��нg�����u�`\[�� E�L8��"����s�QҮ+$ObO�H�f��F� ����6l�xPq���5d\�X�̔�)�.o n0�=+wM�x;���ry��U�ي7�c�E�c�Sɢ c���/u{*����Z!eSL��2�Y,.4C*�9�o��NUd��/V,��ED��O�q��G;�Ϝy�sԷ��B��7��z�;[�
�,e"�)�Ӝ�4 ��E���u�2����(��h⮥X�M�y�}f�`���6L�H�gV����!��^pD��R��#K��ۯ�|��f@E����旡+�v�~~��g��پ�/p�"o��������b؈�ף`���	��	�rimA�,�:
��z��P���`�9�G50�~�m���Lr����h�~�٧��pċ��=�#P�y���hw0�^�X~�Eu��H�kU�=��Qi=����Q����G����5!e�&�x=��	�uj�����`��ד�+�j�wxm�����uPzi�o�8yaB��z��,O�O5KX��O��*؜��Gb"g�@�v�-f��>���q�o�~��K��G�J�~�}b'C�Z[�P������9&A^н��V ���4�v��/ԃ�Hܭ�J^wF&J��1�!�n~�H��U�'���x�b͇-��-�ϥf��S��w�^�E-���#��e���,U��Hܸt_���5J��L�Zj'K�$�7��<�l��X��8�i����=X��8���)��QY��:��H���)vՇB���lQ��Ejv��Տ�m挕QU+"��z��FK�NFa������po���$�F�/|�a���/"��E7�SoR� �V���X
�F�f��$�oC\U�<C�3����
�b�]C,�%�l���)�H�Zɍ�x��Ez!��7�c�� 8�#f���]�D-l��*�|��ٱ�c�%���k��?��\1z�m��*��+S� ��XLN�^��ͽ\/z�p�~*�8��ђ]3y*2H���`�L�ۯ�]��[�)��n��v!,qu΍c�H�F�Y'&u�y�S�wq����բ|F��s�ᾤ$� `�x��9Kt�����Y��/������N�=�X��s�'����8.�7� \��8���{1 >^�M�~0��,�:��&ȴ��ڳe;�V�K�}�[Rmx!1�(05�O�Ev��j�����I�5�+kp����U}�ޣe;�J�B!��Y0u�Wc�S��<��ƶE3B�н_�/
�6¬� �g���o���98���+=/U��`�z�'�����NzFl�@"��~\?S_[��)�5�%���7H�G�2c9�C�JͶ�t�D��$+^I|����\W�{V�z}��
j2����O�'b9|�iy���F�;�{���$��̓>d�DfB����#@�ج~5�M�o�"2�n���]La�I��Oט
`�L����pa,梞B��==�.6�$�@rp�E�E�k�Pȥ�c��펏�ګ�x��MÔpͺ�I���[ѻ8� �#�I�5�l Ų��Ose�d�ۚ,��&	���G����i�ud��_��Ag'̽�~Wːc� FRI�!�tBd�!Pΐ"Ǒ���iӪ� s��X����7�7z}���dӧ��8+�5a�c�^�E=i�������A3b�!�yHJ���9�����W�Z��'4m�>���)L���$��� ���e�����ղ\Xw�ՠV?�
6� T��OWM����_����a�3��İ �+Z�Yů5�#t+|�zw3-�^�	�X�Ln��e�����-�
�h\z�{��Y��6�9��F">r\
�"����Y^�G��d=�6OT|�Mʆ�*p.u���v��e��z(R\"X�rE��^q�Ƌ���?I^,v���_����|?���\�(k����>*G{��'��i@;�/�ҿ�*p��Ѱ�^�߹�]��	�����	���	�=��"���������P\���}a��(t%E��׸o���F&z{�Zp O��P��_!��g�u��\���Duv�龜��1��X�����,�ۄ+�2�Uf�h3��[�+�md��?"W(,��aܿ�ۼ.P�"�L.�ǂ*X�K%��p��Y��BIU���\`qMV	j��`&i��q�L�.F3����R:PNd�CJ�ݯ�l��7�Y7D�*�5���<�V��s4U���2X9�X4j
��b
��^�3�X�X�ar��r�������ct�'����(&���ʶ}�����i���V���k�J�
�����G�gg7�dlV�w6���񜻽^qR��O�u=Z�X�X���]&B�T��-k$~�c4���mڢ�ϑ؞�E�e@�89ϻ����_�-,�7E�o�="�� ґ�ʓm�vN�օ�AO��5(lSH�8�@��N�"�8�^W8kM߈����(�Y4�/Yj��N����\�	��]��A� 埤�(E	2����b1Ʈl >*�d��,r ��/�3K�/$���7e`�g�Cr|	���Bv�"���F�P��v�c��hQ�����ȒX U��D��v`�������tmh�bh�1U%���qǊT_�ߖ��nT?��<��)&���������a]�c�ǁ8;	G�?(�Hb�z	��t���P�zh��G6��D�S( �D�X2:p�?�*�������o�&������:L�����n���6�����0�94A�r�UX=�9C2�pTl��F�	楓�!!BM�-���/������x란7�>yb8ɪ���;�<b��.s{���!��_�M/b�`/-�E�����t��G@Y�n��I����y��&�hT�� -��1��^GM,�7��{��Q�vu7(��u5�|N��84��j!�jA�6Ƌ0�L�*'�0��F��nIM����A=�����DH`sLד��)و.�x��P%���,'�@a��؅_[�����죖�:$��!YgY��Vb��i�R�3m�hu�<u/�
k��3#:��}�Dw;�η��O��M%�Ѩ)�>��~���'B)����9�D¼R�P��\	t�i4j/�3��Bk9�"*V���C�,#�*�9�g�V"�IF��Dq	}�S��	�1@�ܼK ���.MȖt���r�ؽ]�&is�ɦ�d%W��-��#6�À`48@1j�OH���>b��i�z�2�HO'�!u��+H<3,�{5�~?Cl����"�r}�1 �G�r�>�G�u#�}(�KtM���J���8�/���`1��a����mGG�jH#�:H�������q�:O}�Ļ�q`�v*e
L��'�!����W� ��3·:Q�����خ�X�~;���A�8�g��>�K_<�ٰ=�������iC�!��w�JBd�U���0D尚5�z�P��.hY&U��-�U�_$��v��2k�X���A��ټ�QtG:���dh�$ 90�S=�R�5	�l�>+��^��1\h-�ߘ�q�,VQ��kHH,d�����M�J�$����);?3����ƀ�.��}��.fE:�棨b���@i<��f��"CW<=?�ch���N�+Y��\��x�0K91�{����|�i��W��go!��w�6c��-�-�p���o��!�db������F)P���`��;8�G��@ղ�3R�y���RH3(3�ļ�L���L	����}���P���ض��R9�������ݰ��M�
ޗU,�)՝����N�o�O�>5�	�o�>0CS��J:�v5�K�L���p�>��dy�Y�5�(H�@�JL��ڞ����b~Bb`��b.6��PaV�RoV���/K�y1X�x��%m��s,�~7��51��(��d���"9e�ep3~�4�n�Hk?5ͱ<R�6���n$@u��,ZA�r�H�[�]~������<�2*f��ƿ�|����{�RTw
Wm�NO�n���9��V9U�2j!�na�����'I�h, b/lt�Q��`�"��G����v�ݣg�L~�῵u�y/�ATiz�o�
�$��aP6�(�˶c�[�Sgs]�-��+]�%�T	 ���NXn��hz�"	e$�5�X��|�8i�������)Lώ�^�rf�-a����0>�V¥�tcIpsŔRK��E6�R���A��Zj��c�@�o5�O���4��9Ք+�OLB�F��J}�<*	t����ޘ�hT�����FJ��S���Ɗ׾qyN?���j˸��.�ʖ��+�燾+}�t�
S�"p�h�6�h"�D݀+¶�A�ˑ�>D��%)����:p��;�C�q{�:�*�/l�ص)�e��""���~(��}�<�u��4h�ܮ��Q+ ��H��^O�/	Lb��\%�ha�>�1���S�d�������
l���Xt��x�=+�G���]?l��aC�%����RQh�ON�����=Ni>.-F�KX�T��[��b"-��0�����d����a0C�f�� ���&9jM�慊�b���0bf�#d�X�E���tj�#S��f�Ѿ�6Ǻu��7��Y�m]Bŝ��m��h&�;<��y�����Ygo(��|�?��
Gi�&��Vd�uR�>�W�j���OL��ܩhaI\���?fNM����|=M{} 9���*�'�t2�3�Jop_��?2e�)���g�p�4���#���i<���Z'f_8�|f�5�;�a=~j�(�mBS����Q��E5jA�na6�*9���L=��r���!Kx�^G�����2q� �Ѫn�ox�����W ��Gf�n%�ҏ/�D�8���8�1c3���̣���{��Ї2�5�)�?J���!�mOOI�#�!.�[''���j�8+�G��C=dxC(ق�'���@��˃�j���"WZV~��s���ßY�j�R�&A~DRW��Ŵ�������t����H'u%�wX�:N^	��ھn�ʾ~��_� '��sY��J��T�E^��@N!���s>h�����J��= ���R'�'�(BV��
ؠBm���[��5��m���;M.)����PL� � �`I�ܯbU�����Q�>8[/[��R%QH�q�x<�Gܬ���@��:4V�2��!P�A��Mb4Kr��.>)b� �Wk�x�,�2�hM����$�@�Vzjˮ�h�W��j��B�$<&�8�5�H��f+�玁E}}	t�&�DnH��C�Xu�j�<���LIߋ\S��G�P�4��S�r������E�Hg��rqn�"ϱ�O�4�&���u�*C������1!�Ӥ�l�����Rүb���y�4�B�hɌ���mx#\|C_FG� Z�Be#�8��Ol!p���Ԓ�6N�2�6��>ع/�������:e�T���ɅR���ht�(�w�Q_��qN
�a�f6qP�{���̋��T��7�x���q�%{����ec��E��+̎�[͚��eG��w_�/�xn�Z�b��_pق� _�����ahI�P�ō�K1�=�q�l�7�F ��3#� b����7=�>����V�pU��� �ٝrS��T-~�&�Cx̑L���8�k��Y�*���,#������B�
����&�쏵4s��:�
c�Kǎ�D�#~��uJ�6���8�j�^Fw��@	Ֆ�3=��M%�>���n������o��9,lL�.��fRʌ�=�Ó+�`Ƕ=�e�<$��*a����P)i��oq�|�;����֦6/��z+4�d���k�P��Q��:�J�o�*����P�'Y���쭢5�=oG��F*%�g&7}D�(�
Df����(��;�i��>�+�a��[`Ev�P}�������f�#��a�J7W'�o;����+��6+w�ƫ��O�0|��&v!(E]�j�V�X~�	4I+7�~��}�i��3�ld�%�D9���Y%�ԅ�E�AO��
Z#޿�,IR8�
 �w
s7���s��{pw1�F��v�f���b��M������=��aM�% ]�V!���hc�kA��i�s)�!���~v��VZ��<��\�ۋ�n����!�:�w����?�#�zQ^V�k��p@hFU�+]ݔ~%l���o1[��@���ѫ7��i�:������J��v���됕=}f�uG�D3�]�
ꭲ��Gc����8�~XaҖ����F�?Q>�n.��IRDEJ��j�t�a�E�K%}���?�*u=�GO%i�sC����u�U���꽙i�Yэ�tO�������NjB�:7�߃X�܃|�8�8�άki��֖�}nO(A�r�ˆ�;��f��9��6�6[���2��� l�R�gۖg^/R7`u#�^�z Rd���CBe�&u��];#Z7�w���i(�Ex{"ޭ��S���}����V�/� �1`��1�&T,�b�������y3qL8�4mk��Uqr%{�v��� ��S�uy���,gV:�V>ҭ�V��/�9Q���:T@�<�W|��
I����H���ˁ-�����Ε�>9���n_��(�8�E��/Q?4ruTLP+��7�p����(�3�m�R+
�J>ڑF��/  ��J�"d!�ǈɰRG�-�"�:�-�"_���e6Z��vw��w��C�ͧ䚟��ϼ�`�V�����:�A��LV���*��� D"�������x<na�n��,�Cj�mK��u=�N���bk[�=!8J��G �"~
�S/ŀ�g���W'4�u<t�X��Dl��*W���}����(�CL T�Ў�J^0 �>�Ѿ��e+B��k��Q����K%�������^�dݝ6[U��L%dT���)
`f�i� 䲼�u�,�\\]k{ <�%����0H����$���:�ip�s��&Xf*u�qQ�#L�g�[~�ט*3TO��1����2����v-�|U{#����,��H`�2e^��2c�XdV�s۸����IĤ���xZ���}�95��W��&h� �۴�n�G&Ez�>$�bЖ�,�j��z��R��kv,SI_q[|2�=�m=~��j *?�$��kyD�ىO�����9�G��9\�U_F��)�A�ʅ3���}М���p�Y_D����y���i��Ԗ3p�=�?��,c�hdÂ����b�Ƈ�;=���L�k�ɦ�P����]���g��:R6�9n�#��r%�U��Y�7f�M��D>|�ը4]	G��ZW�9oS���})����C$�MW�4 5a���L���c�$� G�?m�Ӄ�y��i�V�~K�kr7X��9�S��=ݠ1ϱ��>-��r��e��fZCS�"���bޒ�|�8�.�2��HUe��,m�2�{hd�$^�*���l(	I�#��H�16i���� Ο���d䧵����ȏ�~�ˤ�u7.\)��bH_��@�l�oȨZ6o<�j*`�s��ykI�DH�l^M,�8g�L<�ҽ�GUVq�J��p�$�r櫦F��j�#�E����,�P^�6��l<e�9ܖ�ݮ'������}�T-���M�����0��� Ԉv+xV��솕4��|`��ގ|��t
�>��}�}���By!�/���+�CքE��>��2B�mܠg\�R���@��%��Y��!�ˇU��i.�����z4rԛ�&�ftP����~=ٺ�KeP�@�ZG&[]�����p	}2�lh���N8F�M��P
�t��������.�i��!r,(���#� w�:�Ϝ��P����w� �Y� v�6NUչ-��xb�_$����-�c���
��IQ^��<e�|ѻ�1sI��h!�-���}~������B����@̓�	�{^Rj�����{��y���7���k��S��#|7��~���_s�Xآ*����ɏ��~y�����mԭ���������b�&nl�dh��u"^[%E�g~o��sS�&�/T���P;�1�����=�B����և�pk �� Qg���
 �����˭œ��T��T}�R���s>}wƭ�J��%��h�R���:�J��z�l�΂�X�ig�τ�����H~o+��p*̘8H��ʑ�#b�_��3�v�ýxh�L��"�m���5�,�d=8�a�z���T�C1�w�����T�cX?خ/�
����ڐ�;$z6^��0�Ƿ'�#%y9KN�Gq�k��ߣ$�fBW�Nؽ�{�
�؇�}��,д�Rʍd�ml3]�
z�����U�����q�;@`�a�Ug#a��d�����L��Գ8,g6؍����}���6�.h0�|������%��.�$��/��o��K�S��j�K����aq���҅pR��C[��WqgBކ�]Z�֌� xv�*��7i �*yiԿPk����Lp����S�_�Q��x��i`;�f��tH�s�5�hW��>���)��ߦ��g�tխ�ܹKL��~Aǒ���{�mܗ�?~��Ev!��c\�3]ⱪ\��֮��9������2T`��2� ���è�u�{"��>�dŒ��<��n��5Hj!rkl�Ċ����;~𷆉������u����֎�T����M�PI�e��V^��mn��OgZ8�*��EiV`Q~��b|F�dw��n�]�*�ٖ/"N�"(8푗7{�Vc��1���ĶY�`��ƾ5�w �f t�u�F<�G�RP����v�W�_��~�e�J�����j�h�*�x�2q�>������t�隋7	dz������p*'px���u�<�/��X���)A�Z�Ymy{���j}L���`LG���*�*�7疔Uf�V�����dY�V9a���7�mAr��ě�黝�n>�/���q��2{�{��Цҳ��].���y�RJ�8W���Cz�����ց�J𵐗�}I/uZ��=�DpI[��xr�a1��0�K�/�o���A����?2R�0fK�˱N2+��i��(�h��8���3s����&��l����dpI�ᏃOk��k�@�M[�;��&��oʋ�k���zV��o��w��+{	'�5�h��a��!�����40�D�z�q&(��қ���(�>��v+X�wnK(�n�`���h�"ή_�\R��v�-��T,���(Cց*5�E��"�q��â��$P����ȶ��z�+�BR) b�Jҿo����@�(���2�[����}���N�J,:L"��&#�WjE���t��zj%J#
�TK��|�I��K3SƋ���N����k� ��Ř��ƍ'?�0���g)u�ev�C7D���h�	*�����h��߈!�V���~/��D$��0y��iKJ�th����=�&p�,K~���E�޼�hۯ�^�vk�5��~�^��<zr�bZ�y��J2�Lҋ��%�>scK��ϡ �����]�Q\*�g?��x�hB��g�:A�8OTS�l���Q�7�]���9h�A�k=j�?�)�#���+��dU�Ġá�WA�h!y��j��zB�}X�=rv�1%���p���Dc5��������*�*&o~(���n���[ɛh�3_���E��K{��Un��}J���)u�y�1�R��6��"?1+ů��6$~$����I�n=R�4��"��](1C�D�ѡ/Xj֯� �9 ��Y��v�������Q�1Y�wWi1�Z��?�j>[�R�S�����M��9�V�Ԥ�ِ3˴0��?�t��VIN���	�h%G��<���l�~4,�w./��g�ԦO�@�sf��%D�3�C�R�����t��<�Z-m���\>USc�q$�R��3������Ҽ�$G5p���EB�+�Z�-] �Ϥ����}����g3Z�U������1%c�L��W�hA�X�������Pȹ(Gt5�V\9gS�������v���E��5\�2�n�r�#*�Kx�s*^;�_�uYp�n&�p��`��G5�)����6�Ke��8-�J��YJM��?<_H;���,֜����@r���~~#�"����<YӮO��O)H+��N��)w0W��Y�+�^��Ǳ	y'7��L>5Q�-�'}�Kw��<_|l����\���7�I;#�v�t���,9c�2�����!.���S�!԰����҃'�D�Q�OoӜI�W]W�frhL�~�H��B��}�P˷$]�*Z�+���wn��� �!Uv�3�T�ΐ8$AW_i2nw�
S���W&�J��m�"��!5PL���@M6E�^�t�ϖǈ��L:<����QN�3�U{;�x��X]"��E�<K�7�Î-ԡY�ƐߐC'��W�WA��ǜ"=0.��K���P�<D���'s���^�^V��pv�inM;z�[�n���&i���	�����Q����2�Xܥ��@}��뮵A!9t<���Їy�U1\]��{�Orͥج�B&H]s4+VC�vC�aۺ�,�H[| ���	��{\�mX�J:^WJA0d��|�+v���1P#s}K�s�̻��z������.�7�!IW>��om�ڪ�5Ȩ��(��ԁBO礮�g
u�d��,>����sܑ&���dh�l^!�D]ɕ�� 1(m�m�o(����s��5H��^ZވH
vų��|�L-���ܓO
��z/l��tZ��<��?���l�$x���=���~�ﺷ���aʘ�, ���+n :r�	%�Ve�4f-ѿ@��+��F�S��.!�4�Q�:�Z�
>	�����]~�NV��n�{_;��cw��t�*�~����+��?��O�]U�RB�OȖEߑ�?mA�^>�>vz^�F�����m�"�@���f�2�Q�d��{�x.�� � ���� �)��������\��m	�����ҽ!�Q4�+�fؒ�K�;1�!:�أ��_B�0<���@��wI�>E��;|Ϝo1Ĥ���q����֏�S�17[(���kuO�!�Tۄ�ng!��c�bPqe0o	D2W�f�R�u�`G�6�֙^`�\\]����y�k�zN���hV�I����d������qFԆ0�C�I�K�l���}{5������h����^|�qJW�>�����$qN��"�20���t	/0���� ��F�Q������O�(lE���ۏؓv��7|��9.e�b�ik#�&t��E(;@�f�9��nِ��ċ��>�4�<S�r�Z�/�`A�!��&9���ƨ���En���1�M/�K,��������0�_�4k��y�|)~`|��o�􏸌No�aL��)H:�8!���E��nJ�8l��P�s!�u}bR�XTߛ�`V|����Z��$19�N�MIc�K�ՒiH��N�%{EZ��@�����huT�����idO��NՎ��ZS"�n�7ǋ���!�Q,GD������h���i/	�nx}��j��v2�f�Iw"2��'�i�C�y��i��]��D~3�o �"��L��Xk����3��
�X�Y�7NIE0
��y<|4w���%)��Z��G��.��Zug����Z�DD��h�P���Fe���E��c;�<R����6�jo�����7h����5w�tZ�z�Ny��VI8,t��$���� k�x9��s�)MҸ���3vzz�[U���~�E��� ���o���dĒ`b�AN���>(�9h��R�2W�jR �$�e��U���0�|��7zr�+d�*���2,�YK������wU密|R��+�Oŕ�W�ӽ{�!1H�8iݩ�KJ��n+�EY���B�	MRضDx��4�9�L+�"#VD��X8�9`V�*"61Qb��ǃ������<tP��9y�"��b@��S��*�4v�\�l���=�,\[��]�:����Ȓ���`N�l��m�>F�W�z�)��1'�Jta�9v C��w�Lf���E%�OA�0g�(�%ge�47��ʾ�\A�D�1�yAcD������=������i�}�$�
��	EC޹������S��~�G��p���L��j��6`�Pь�}�"�����*�+�`p�w�1���>�o�C�'��s�h� ���xF2�����{��k��O�%�N��v'�#V�rh����v����}� ��ٶ�/�p����.�K� �K����3���C�:\�lA�.�/�R�xUk�<��3'.r���@���H!E�,������=�2��|]O�F�h�]G��ȇxj�N^eX.�%LXH�A�����8z� �6i����U�n
�vׯ�Itm�r��bL��_���}�����Hw�*�0�#��ӹ�!ɹD0�`��=���@�i�6Z��
�^�D>��
}���ʋ�l�R����ɲR��g�v�,�Ы����bU���5i���t�:l�+�GRQ�A;<sGK�i�@0N1���/ͬ�d�u�3�>IRs��ӂ¢u(fc#��-MY��y�x���z��Q��ge�_��1v�B��^oV��ڞ~�ʼB�5���	���S�zl�4@ҽ@��Y:��&Q�S}���q�f݉�KMG���ikC���F�*�h��K�ǝݢ�?r���{�z߲�}-�
`���eA�z���ʐn�/�ֻ��!�P�=`Y���39�}v��֢�
!�P,�T,��É��g�_3l�f��10�x���,W9��&ʁ�=��x��p8,E����֢���P����j�	�M�᳏WmԴ"�}MÀ�O]�[��	OG� ���0K l�4>����tr�"|����'�&?�x���
�ٺ�v�hv��r-��S��\�𼳩��ʎA������R�0[��K�>�ZI��:����9��߂w�QƖ���g#��IO����Npr���z���fʻ�Ƞ�I��F�f���4�k'R�e���!x`<�;j��d��r5�3��J�V�x[Xɟ���>'�4��~r��<�s��a*��r�BD��!H|�1Zic�^Ѧ�Z�c���G_�r&�SX��$K\2��s�V�3��m܂�2�ss�k_��>+��:�A��mX��Ѿ�������1�Z�q w&`;S?������tB��G����� {���d�c!������(�z�`���/��G�rQ�'l��1��Â�z���7iq'�qvԠ�"�+U����C�~˞2��VB�x �A�
�18�ei=�|b�~�!�t���Vֶ�:I�m�$��?���t��5���3�� �1^o���MN���~�����}T鹠�b��|�4L�1IV� 4&�0K�b�ҡl�nձ{����;wS�S!�*�Vo�Vs�ۤ��?��ݕ� �d`�c�An]oΘV�R��t�ھ�~㰮@cķ��VԖl�m�E��"��I!������/���v3hA�,���p�5b��ޭ�����]׬(k���9ݏ5:b��{����� ��&s����j��h��^	��G�>'���:uF�K�}��y%�18���]�I��#5~-u�y�6IE���S��hO&���PgML�x������͞�Z&)/Q�ܲ����\�/vw����� �@���A�@y�Fx�n�m����'��m:�p�ϭ6������YH=}�4��y��a�Y���_�_kQ[j�|��SY-N)Գo�0�ړ�u;^�;���3:`�[�L����c4��Mj5��ah>�p����Hb�� �E���zIϋ��=��3�=��վ>�E��g���C��r�g�G%o5�m�y�_���t��ͷ:_6�Ђ�ҡ�U]��� �0M
��1�g�����	׾�4C��j]��r�K�^���N��/Y�]2��.h�=��>0n��68f5�A��`��AOhՃ��͎%\��km���hi#W���ԃ�Bjn��]H�?\������80y0Ə�p��?�#M�o���@��V�?�V��P%���L��n���RBo�Xv7~}	�%k�c&�rf����c��T�¢��h��p�du�,;+gz�RL�<�|��{�8�X�?�n�o:�݊Ӳ��մ��!n*�)��@���-T����	V͈�n/Au���5�.bн�/�i߸N�@��3��0�G <�)�&z��Jz�I�@�$
%+�<��-���#�wpO��̸����Y̟�}�6�:ۊ9t_8�n�|u4����Ż�ϳYj�� �5���d;�PpkS�ܵ���	^.���Ph����d
0�n�"�X�OwN��7�9�������CsUtSLC����hk�'����'֯�������OEs�MX�?J��z�'��۽A�D�J�Q�����a�KO�~��\�CU0��m���x�;�7H�%f��'F{�g<�m�>V�w�/�u��6�<h��n>У��_ܢ�P Mg�'Ӧ���҃�Y7�W� yr�^�Gg=f��\���J��'�2ge�F�r�<�`Y�~���L��=��f���|�_Ϗ@',�^sP5vT�`����wܪJ�����u����MȂ��X?���\ �v�������U�5]dR�w{��������a+%0ܢ@H	׃�Npj���f? ������"�p�5��"����1��l�1�}�Q���~��5��0���I)�c��M͆���D���{"M��'��<QO�Zm�}�F�q��V^]R���C�[��6�pJD�ԗ����"��:���B�h1�6�^|j���O�c�}�ۙ4 �&WM��;�
��t����f����jO��U�,�%&	�2�U��F˿��p=
�����.�Q�����J]�����\���q8q��	j��9�*���Gr�����go��|72i�7�V�f���s��c�cm�D�^/߲����	���Υ�K�����]���,v֢�Ng��ggpA{�~����.=�����6�ц�Qq���jR�?�t ��$���bG��gM<����j ��M�nY���r�x�$�o)�:z��l�qA"�f��x��!뱧�@v�9D�������f0�3��Y�@B�a�Y���)l�׸)��s�3:;���5���3V�>꿑��.��8{�8�Ef�J*���D�J[L�La��~ñ䖞��^����dX"��u�2�̟��sݹb��8������{�,�E6�z��ڮ���+	a0 �3��L����9�����n�� 5�|��P�wB=Lj쪳tc����ӷ��.�Qة.�qY�w6u��)I�2��(J'i��]�[KO�����Ć��E���,��YBm��g3������cA�g[̱W���ɏ@� ��G�V���M"�a˓�r��̌�2S��#�s5�FF�n�m܊r0��aк����<�5t񺓎{ˊ��X�2������#��&�L�G��).�k\�N��F���
W����k$ٓ�L5�g�@?����89-\c@�M��=7vBX�|���f:Yf��#�+����eu�*Ӟt��X�7,,N���RـmL\.
d�����t�n��[rf"���OM���5�Z�ىޱ�ާ��d�~�ڋ��0>���f�G.�ǌ"��� ���
�~��s�X�<$+ʐ�k`�C6#$��v�?�)���g���Fe����6i`����I:-�#|��L�ˮ�$a�;aϙ�5��8�mC[:�s�yE���0�->7qp(���V��YM�u��v*��S�H$O��6Ss�U:��݌� ��+� 8Sʭ3��?C�*_<��0t,��Ќ�9^/�W�_�A�"b��
WAK
�ky�'�޽��o�?I�Ar�zY.F��IC(���b��0cǪ�Z3p(��_VTqR�8,�"Ȏ�[����9W�$��1�5���_��$Krtkd� vz�J�j�X��ٗ[_Duk���(��b��6[�����B'���mK	�W	Я�$Z!OKrN�����#��[�2���X]���{�pU��}ص�K5�i/:c��d��� �$=��v����i�X�;}'d�ZU��3�dK�F�}P���3��&Z%���;U'�6{����X�⠄}��bi���CI���l��6S`5��o��s��Z����ҩ��[�jק--�UV�����)1��W�����:��ԊE�l)219jUh"5��z��y��r�E�0��=I��������
YD[�{3&�Ȯ����߳�m�;��]\�nJ�tW�O���ՑM�Ǆ{I#k��B5��v'>�C({j>FwV#8N���_�C��"7%~�OL�
�,��@"s�JRHb!j�B&��[>I��L?Z!�@�9[�=d�;V�00�/3�z��u��Ǎ���h��ߵO������n\��*��R^F����̳��~e*FǓ�(V)�y�M��nd�T�X�o["\�O
e�_�kG3��|�jG��Ţi�?��⧻���Y�G��,��qB�m��PF@�A�K�Y
���=F�@��4>WEݿ�ц��Ek��j3̶��9����F���F�� �U�/�"���|���Gm�u�W�������.��u)��f�{o�1��
�0L�����p�Y�dU�K4�s\�̻!$Hb��Â���f����[>�_�B���nh5�SW�HO���l	-��p�h=0�F5�M�FW���f���W����MȆL��j@��\tkD�J�G"�ʨ���A&��%)�u���yh|��������u�$7zk���1�Zld����
����[��>��B�"K�!;!:��^:�u��_�b%�8�u��ρ�/��s��P9&l�	3lJ�8�Ԧ]�UZDy깒̃%jIx�k�|
�\E���K����Mp�?=��h"��,�����B��eƂD=��/X�����fR87�y����=GNY��^��U8��ʜs���AD�`�0�� Jk�f�!2�ս�-U4�7�%hE}�%���V��"DfF�2�]G\�� ��RaW�(9/)�.Y�Ѿ�/��6�A�~�mm��j,��5�,�cc3�;�m[���@���?���)�R,ș���Ѹ��4�49}�;ʀ���%�L8��A�+z�-��z��|c�[���%M�!_}�s�;���$�����E��.�. ���P岓گ^d� ~:InC�8�� ��9��u,MŁW|s�k �B/����?��3�,+v=`�GM�U��M��_$5�n�:k81�I�T�@��f,cL���i��q�F��Y�����=���E1�6Wˢ%2+��iɮ�Wp��,��S�D#@�ue�=:��a�Ӯt�l7�CXtq����nd�T5 ��Z��3����q�]@*ט�F/��sMnn��C>U�e����X�M����[�Ǥ�������`O����y ;��ބQ��~�A��9D2DV�f;I��i���u&Ȋ��m�������H`���� �"��_�"���7O���.�m9Ш>_O�8:U���:Xz�X�/�3;��g-1�03��_�D�WД���A]�zG�"�$��@Q�� �g�;��R�+�\����M�-�d딐�-1#��`������ac�� DZ��ia����$ȴnP8ګQ��a&�o���X�~n�6��(�z��)T/s��]�+>B���#�U�ZR��9� �'8��	����GĲ��W�1}��DGr����i�2�#��� ���h;�N6��vp���<�Ɠ��*{���ߎ,�z�=#�|��x��2�������=� ���^��;s����A�YNQ���% �:A�6=d�\|%�B��+d9��	���K>/���ӆ���U$���:U����( O	�!�l����z �h*|��$H+0~ZSH�Zǟ��4�V�G�A<��r⏇s�M.�����w宑3��Lp�t�r���ZA�S���zi�|�e�2�c`�PW�M�#���M�����`۰�y)V��w;��"�����7Qc�n3 ��g[���E��A~'���[z�aJ�Ʌ9�iLxj��Ϝ�3e2v��lh��tB����;�){�QL���3�4
$�N��$*GRT���Q���Sџ��An�5��H�� @��U��=x6��5ߛ��8���
A�	3��em�(,[#e�rB4��-�������K>��!W\����0!���܆�%k��l�����pQ��҄}a�`'����<i��������zs�]���0��EŁHe�'�lR� �;�]̯��)��P��b��mA�#��� 3���Qӵ�����#ͳ��8[�C���j�e��G��zy��Z���Z�W��x�SWt8-̾R���ҿ��a'���-�U�����>�[>R�V� j}���j�.e�&l�Tsݱj.�YY!����n��<2�~��*�ޗ��*:��N�}1A��ʈ���m��^���*Զ�nT:��ԐH]�ĆL\jW�F�o��\��L�M	�K�UD㙅\OU���+|���4s�152���cM3�ΈS���|����덎�1�]���B�X��O�����)nO�/��ue�{��I
57Nd�J�e;1��}Bִ*�x_�Xн�L�m5ɿHt�l���9B����3�>�P3�ď��fǮ�\T�:��l(/( v�8[/�F���x��4ZĈ�
�'{�ʦ!/(^���]�	�y�۲�r��Y�S*˨W:ޒ7�xP/*^�M� 4����|��Ii'Y�oH�ܙ��������3<�Ry?".�E���s�������K1�+���Qt��34_VL��;Y��-�Ou �Ϩ��
��B�m~@�a��KZB�m�DIh'��HE�#�"D����9}���Q\hY�>��d�Ev�;�"��j?����ųWz8�+�fs\���-�����Pzw"�į*�y��7c�%�Z�_�0gW+�%��%Ia��{~D�R��m�iG���f��K6)`��YI�{΂�S���i[w���j�f��1�K8j�N��4lq�kޅ��w
��n�|�Ͱ�BF0��M���(^�0����)G�x�������"�t�@'!��BQ�V3L)#Zj{�<S�7k�r����*;�J2G��[���L�v������:�?���o,�P^�3o䥔blǍu�%VTjD�ϗn�N���%D��%�FӔ}/[MV���	��dh��<k�����Y�e�9�|�p����H���x>�&��\����H���5|�f�V���>���!����U� Y�7@2��8��N��r̷F��g$��H��9�N����x,�N�0y���ֵ��	!�E����1�����ͱc���C�����һZ&Rhd�M������tZA⁑��\�����4���$�W'���ĺO�؈�Li�G���ס!�5��<l�z�7'��p�o���s:qA��IT�q]O��`w������a�S^��Y���7�]�}�g��+>�c�TZy��CJf��}��e������){��deD�P4�l�� "��y@+|8�\���5����=%�-E��iX�U�,/b�o�"` �mڏb�W]9�c걹Fv����=�.��;ʼڽ��^(K)d xG'}���8s݉w�]��m/*��J�����v�<��CLi��6d��˩�x�u��W:2�j�_A�8ѫ��"��4v�F���V-dE�}�Z�MQNvm��u����FJ��g?�o�մi���{=�d%��si��!'���NR�O����
�d:�A�`I���v[������K�]2IO�9��u=~�R�y�Q2pEX�%�O����X
5J�߁ {漩� -�/>�r�~�ܡ;��ZsȀ�ÿ�S X�@m��w��\�#�'z������ġ#/�|���q�Vlh|~TC��u�k�Z%��
g� ���I2`��`a����H;�@���76����ރ,s�T̩�	��M�@��e�/�'^E��(��X��d���=�D\.�w���m?�.���,dfp�m�DK툙:�*�f�d�'��)�W�)���tDH���L���*ˇ=��Xf_{U֬��N��xq��1;1�r�,�B��hz6���)��GB	7���v�'E"4��F�6H��4n
�pZˀ{�)���b�yG�(`�4բ��Ѽ�����m
����o{t�B(���L��_��戋n X�)`��l�����0s 	'ռ��1)^>��*-$������r���D�j7~��{���2ze��iJ����/�>n�C�&K��@ĆG���e�q>Ⅵ�oN&RV+QѾ��8���h��»��2�α��]�,
��j��lf��K4��d�Կ\-�4(�8�\)gM����:�� �{њ����[is�s
���]���)4S�7�(��7��x�b�k�*f�����v�g���bd��.�Ồ���uЎ�av�����X��G=�0�K���-5K�J�0�c]�
�R'��ٸ����m��e���!9C;m~�t{D��3�Q]s�X��f5rRC�f�4WMp"��jZ�%���.ͨuG���y�ND�T���k�@ ��	�ӊ�K�Y�ct�x�r� 6�2��*�#-Zc�����r�'X��0�iA1�^���5ng��T�XPSb� �)y�M��g>Q6O�<O�+=Rqo@�>:�+� �w^�I�]>��k���)gF#�|�$2�ZYH�{Z�!Z7��h�3A��t��;���bB�����	�0N��8��J9��`Ҡ1�8D�)�?:�1J|�����pU4��'x������`6Aǖ�_c�C���s��~ؤ�q]�(^�N��S��b	��,�S�\ػ��ЬMy�Y1�:��B �P�8Gs�<e7��	8�귤��j�PV��!�a�O���*O��:�7V�l�$F6"�&a�
Z�J�}
�v����B�B`��f
G�� c���|�h����Go�ϣ�NA�d�eJ�k/��0}��+S�ic�<�T^q�_��R�%]X��wS�u���G�ÏJt Kŋ���e+V���E������y����v���5��B�T;�E{��I�rWmµ�R�<!Q�_O3���:8��)-�-�ZU�\�{Q�H3�	��|�zQ@�S�u��l%W�υӚ����XT�<�$FO�(��l��6�5+���Ye�w���*Ɉ����R�0��QK�},���woB�O%�%�������P�c����������:�֎�Y'�&N�"��I3O����H:��Y�,_�ɓ�{?�/�R�c�F�I�#����uF����}�Nm�3�ũ,��J�5�Ԃ��U��B�dl!�vPK#o�I�V�`I��&�ޑY�����Y�@O��C�N��N�/}0�D��o�z~�#�?���:hl�ҍ�@�����B����ň�2!�{S����ux���}���������5ÞH�����B��E8S���݊��o�t0�AGf�1.��6[��gB��ÉSٟs�4p�ͯ�W6S˳���������D 4�]���w�r��ME��ڋ�r�Uo;���诏s��te(�@?S��:�X�{�����#�uЕ����k�T��]M���-?��`&�Yk7p�= 0�%o5QH'�8���K��OJs�Ϝ�bH����Jǯ���"��!���`3�̱5gJ�:�}���'�+�[�ݓ
<�#'g��� �`�4Z��!l�O�b���`B�S>jgN�& }Y�nv�Ҫ�'k����
��-�� {�_�؂p����e�7@\����q��d��"��W!�ZA�3ϋ�xbژ�K�{��"K31�{��4�Q<�:�?�(Z֙�"Ǒ�Lll)��-�8)���Y��]�f[�q�~����=�ƛ
�4|Y���]Gʌ�m��'k���U���?i_���B	��%�����7�Fq�F�4��ᦁ�LC� ���7QM+	�E�F>��Vxb
��럢�`Q�X��D5V��I�ل�h�q��d��,�E��m�zI��: 5L�� ��9:�����j���b��]BR�� �*������t��k�/���	T̅�{�
�	ޫ�;+u���B�0-[����Q�Q&�sٛ���QS��h+��ڌC��oC�3,K,8��"f1'R�x��3� �;xQA��Mv4���Y��x�Q?uW����#�V�H����`*r
�#� �q����cwe8�����k�G��o�֬a"��
{C��Tq
z�v8g	8N�r[���$_�&*q0.�'=��������)YqA4�!�,�|���ϐ;!���c[��|q�1o.h
7�",(�ۯz�z�&�:~�5y^�,<�Wq2ǐu�!YvC`>��T��)���ɯ�*ˠ�|����0ȶ�;�(��+�R���T��w�h���;�O��i �h�M%����Oe�ݚl�&ڮJ}�ϖ[��9/Y�EД����:,켨&�P����H��1P�6�<Y����mvh�+?Ԍn�I3UZ��آ�lu'�*ZEGE�#����,����|ؑ"�����/��7�0�
p�%��_{��GECʘ��1c�7���I����Cb}"��v��п����S�O$��
����,�XH�o���){Fٳ+}%Jq�j��yY��_O.
�>�H2�Lo�Ѧp.�/�K2h�|Y
dϋ?{\K����: ѫ^��!0���ݝ�S�y��� y�Td�ws��R]�����?��bL�� ���5 �k�2F� �����p�,br�]�"Z!H�:�s��}c1���F�ӡ�k#kp�-��beKf��G����ߍ����o��4��z�P��,�pP�q\URs]���w�!���h���IٍN1VZ��bg���#�0t�{�S���2\9g�*Q��y�'���p�截v�K�+���Q��E2y`J5i������I�.R��2����֭v�`���_�ŉ�w�n`A�B��WG��}��LQ1�E�
��Y	�9)A���:�l}<�jh�%1[S=����R���0�%EFe,"��+��������Ȫ)�\"W��ݝ�9�=f��x=��>{R<���+b�N9~R-�6w
"M.��`߬r��;��n;	����4�\�Tf��d��.�B&��$�K-��G
a�HOw�|m,^�=_�-3�NQ�H>7[2UÝ���\_�\�����Q ؆�!9��&0����ښ~�.��������^?H��?c�W�&�`���(|� lů�0�Yсe����)F��cH)��=��y������95V_}*z���(d�\���|��N����q�s0�;%����F�^;��̌�tס�C���Fل��gI�5�Sc�5�b����d��ٲPv�f��Cr=��(1��S< N#.L�	Ü��=4�,A�e��;�4���g�4#��Iw^�x~��U�����#�dn�+�m�����4[m)�4v��*C~���AV������TA5���xȄZ���odV��$�"MFƩ����J�SamT�@�h6�w\�y6�IX���QvP�v2��Ky(W-J�F�ݵ!���H=L*�"n�Q�v�o�$�Or}j8R�O����Igw .���7N�q�|��徫���z� ���rX9�"������)�b�A|^N����ф"�7I��bb�З�i�w �=|P?�@(��J@�'L�H5�h���p�>�G����Җ���c�/u�Qja����Z��N&�V3��a��������!�ǈ?��s~��B�dk0�-�PX7���P&�jxer��~�PT�!�/�W���z�H
���1Ve�_a��c`����K�=. ��뿆�|�i��se��CiO��zړ��~��{�~��6�[�� �<�ڄv�`�Qf� �%y#�1�4�xwG�(���yc�Dhi��4�[�8|s���c��;.��Z�� *c2�V�q��3�U���׬����*�\��c}ʑD�T\˱��&\e��V��+U��a%lBwa� ��n!��O�^�c��֐��2^��� #�����-��S�� �OE7[�,�,�$�;Sx�a��K�/e<9���p!l��һqh��MLW==���+p��tÚ2�uci^�:Yڞ����n>|&�C4"�����=fȪpZ����Q�_3�s�l;p1��o�0�����N�#M�jq]�������T#��bR� ��H�v�9�)Se���#Yh�<�)�6[C���: �ߨ�v����������� C|�#..h�B6ft��ڃ�X�?7?b iFjT�<�Krdk6|̂hj�5��`�nMGIx0	�.�}I�G��%pr��Q�D�`'���س�6�i����1*O�<�hC41�X��ll��͉��K�Ж�P��.A����6}Â��>HhgV�P���J�z�񲐘�T�[	����v����.���J7� �}�&�;(WT��в��x hX��(%+j!���������9�B.=J5&x8�UR��MjZ�T�c�1o(���n���1��5l7�^�9e��1g������4�2��M��|�3&��S�LŪM��^>@��^���d%���W#`�p�r��[N�����4͂�H�.�9� U��eL��k5d�\A71����Q����7��P�w+�d�d���IE-��M��R:c��6�@�%R�d%GT�y��:���m��̏H��N��e�:�B�k�!�2���I|���ok�̌0N�e�n8��t8|ݴ� !}����)@м��ϓ��/��ā<��؟�op :�1��
NM%S�$^N�,��.j��BꝒ�A���cT_z���y�e.C��v�����#���}O4 ���6��7��#��E��'i�k�an�SwM5d|�j�2�xO�p��֩s��o�p9 +0��D�+��Y�T4`�/�!�Y� 	̑	�`f
��G]�A��H��>��{����3j�f����$�Az1)y-�<p����!.!�{��]o<}�2m��ﾛ��ŞB^zt&�,8��v��kgd��\\\��59��E�Y-��GÒ�#պ�$� ��D��y}��|��a���_:�� n�"`7r�;�`�TfpY��X1(����<�(�c��T�SiD����w�k�Q g��<�\*u�9����4��8_�H��R�9��M��A��Uݕ�~�n�l0��OŤu��Ź��46���B���ghخ�Wǹ9PI�$��&d��L��r�'�/pĵ�=�EZ�9�rl����xwhe����k�����Sh��,��&�u�k�V��U;�B�[@�6�S�.k"/���`�tG`�5�]3�w3]��� �� =L�t��C�)���_L�7����A���Xd{k�4��e�X�3����t�M����7��c���{5C�xt1C���7��?���y�	5�L��bKݨ/�gC9$(�J�o���܆�y�O4��G�3�HVv �wl�D
�����?КC�z:�
��3OG-!�+m�:a�R&�w^P#�N��D���܂��o8Pt5�߿�$�,{�O���+Z�^���ʣQwU��1j��P�e"�bS�h�h�
�8n�Pw�?K�k.��5F[U�h{�Cx�s+|����.!f��g�nǔ�g���U�?���,�N?�mO	�0:"p1j�jT�ȃ��/Y�Z�~ټ��i��uc���?��%�Z���X�iDA����5S�Z�Ge�\ʺZ}�/��os�K��a�r>�x��E��{|A�Tkϖ��C'�|Ջ��p��t��{�c�$��7���k=00�@��b4c��h:����!M�G�`irz��r�D:��xK����k���t�L���1�T�|���dX�X�=2Ef��Q�; ��AP��orN���C��"�:_������,@��ߗ�)����*tq[~M�<��p.�0`L']�{H��iX�Vm$ ��u�^��P<&��Y]������Q�m�#�F�}��xk8t��@����ZhB��zg�����|�ΚJc��:Ҁ'Dk��\��o8��jJ��S^�}��MG�\��~�1�	�꿴1Ζ"����p�=-��D�:~��{K�MA��|"S�_fQ���l+����9l�r�����Nm�������t+�j��F�n����9�\ġ/3�nH ��T� 6��j`ò�"�U��x����]"�VJ�g��Qw���4���D˙���4�8>J��2_�E�s07$z�l���� W�e�_j��C�JTK+"WncH�3���/@���M[>�`9��|^�(C,� �.f/唨"5U�]Vօ�A_����R���U��}f!xI�8�����"u�`�\K��V��� �]>
F���?�Q�9ʐ!�lpo,�K�d���55�	`[����-�9�����_�F>q��;���1�lKn\��дL7&!��5"D������{����Iy�~��G��~x�	�tjKA�a�'�L�5�W�O@Ǒf��J��e0����
\Uw�х�]Q��(�+K�
�wx~�I-:.�	O$!w�^�ګ��ݱ� e��	���UD��Q��),���M�z�)�zR)�4Kbe~l��`������|�8�ܳ;���":����WQԢ��~��@ye��Ug�l�`
U�T ��^����^3P}@�B�pux	怲7#˥yA\�i0��dS�a��k����j�2�a�G2�u~��-����G������V������]��>;_��] � �/���Lg|�`ey[5���n�
�*�UX�t��)M)��T�����۠4�F:��p?�'I܎��x���<J��������̟���~6��EQ
Z�:�	e�?>L�E�)�%mlWD='��(��m(�%�ȅ^���Қ���k�I`�TWMS��&{�	�P�#�g�2�U3w(z5��ш���cЍf�e ��t���'��+=$�B�R'2���~>h!�W��爧���~B���zD�;�⿪i�����/����Ȍ�:�/�n@���S�:���N�FR=0�gj[*2>/L���*#��1<�t�[�*L���mEo_
��`���Q�d� Q��,���D6
��2q*�*'ǃ1�;�)&�Cu	C߿�J���m��%��O(Y`�<a'���*O�;=�!�O�]��Vٿ��Quw�j�T��3��(y����3��e�o��8��9����e�5�8q����a�5C43�Z,/�ޅ*zv �pbB�
E<���N���pz��=Am_B�%�h!���ԹSS��޳�)���%�ۍ�u���ۧ�|�$1�"2�����]������W�ѡ
�Щ�S��%�]�Iȗ[6>b���%�<Nq�B�mn�������N&� �i������+xzy��3)F>���� �%��c�-b;�9��i�:;�{��l/Ǿ׎���&�Dм�[jmEC��`��
+���+3��ԛ��1�ݶ�DRBt������F�F�Y!�Q�S��|M���'n2��.���Cw�r��\���}��ߪ(ظQR2�=$䣅T~�{��A�[<AK:��s��͝q�<a�k�x�HcVU�-�<U��jmz�EeS�0K�ʅD%rc�l4��D֙��������y���˳͛Ӟ(��6?I��"q"^��k��s߫N��8m$Eai�ٌ�����$��(�b�!�:+C\J�Wn1��[��ՊH��Qv��R2�)#�@����%�޳�0�7_㢵^@o�|m/� V@���|��8��@�t����^�{�.=�;rr�����f��&�_������ֻ�)�M0�16G��8~p�m���]��֞_���c��5��0o'Y�lI�9b,&���Ql��Z�=�x���،5ų�@�x	S��Δa�{���N�滈��7���4��BBr$` 9��-"b�%���j���|fn�KIE.Yuť���7��{OD�7��"�vھ���Ś�;�u���݀-hB�k�d�ԋǔ��qh=H5H^�|�ڌ��低a��;�	U�p������"���d"A�N^+%�Uw!h�$�����>�l0|�@�$/np��p�1
ꎃU�Y��[K�/0n��i�gvd���2�W��Aoa�W6�a4�+Xu�Hr	r3��8`կ�x5U����_��`W.�Rzě�r0Z�$`r�8�dm�k�p|N쥇�_�"��Q��c�Ʋ�W�>
�H�/7oh��@V{��O|ى�����u�5�H�Fٖ����!D�ǟ��"���LI*`�y�x`�ĩ>t={C)�	�3�ը=A�W����:lswy3�I�!Y;T�/"���5e��I��F:��#�e�g�O�"ʋ��뱜T�huXg��k
%�5M�@"�t���H^����J��� XUp9������M�q����eV��?hs�e�l����\j��#Q�3�!~�e��u�������L㮳o����+QS������!}��S4D���^�>�nӤ��Y���ڇ��$�$�nh�s�4����@��8TI���a��!iX$"B�}D]:h1r뿓	����x��6�wG�\�o�����x��;�vwT~��k�d�9���&s�lE��&kp�Fߪ���Si^�� ��-G��}Y4�tɂW\3�Ovż �	���~�E�b�1��y}#��;]���X+��&��Xt5{��+�d�&����|��.����h�{�|�\!j��>{Vݘ0B7�]X%�ӁV�� �X�0Uj�.!R����O���.���D�Z��ܗG���7�O��(1'�Ă�	wT���^F0��ʤ$��[���u!�I�4N�t������|����oO�N���jɚ�SG;J����<0�~�cKr���SŝR��q~[��|��=W>�Rc!�ܺ� �Q�L~��� %]�~�[�,���Ov �T_��Q��Ri1%��*C�Y�ӫ:d%\Ѫi�C8�[�+� ������o�������#�9�s�����-�L��u#�_t�Z� �{�p�=p<���m2�%(�n�(O<�S��9"�ӕ��T����b��\ M��d��;���og�Qn��'Cc��(O��_yV����y	.5�Y&y�Ĉ��7�LVY|�^њ�ɏZ�����}�X[ۜ~�)�V�����n���B�<��D=����
�u�l����z���ko��T���te�S�V2����ʩ~����~ [��*�o�s�c ^�_C\E�?ך6��Ԅ��S�'��u�!��ڝ��z�LD�7M��w$�X,��X��p|n�'gFr��;&nl�9s
��:�w� �*g}a��$�����d�?��~�N��8ohh`e��F���|3����3
U.oG����o���B�I�Pw*cZ*xt{nw��9�h��������3��uB��v��P��Ј_'$cS��o!�xe'����������Q���Y���Y��c8�f��pfԠ\5��N��x�I!9��ʨ'x���F٫��f�0���?'-�q1=��d?AL���%�n��0-�<ע1e�����(����v�
8�c��r��)�M�x�R�B̠�� s��&������m�1�NBwZ&P�6l'�V��TU� &}:�{<��#H���@\h��X#�G��@�G�L/�Ew�2!�C.ގ���k�X>�2�n4��Ab��95�T0��+p8��L����9�)ט�)��a�\��J;Y���Ѳ�Q��^��ߟc@�Nf��Fr�������$PM����ڻ5R�O��.Եsouq�5s�@��6U�4��T!�@�b�R�Ո՝:"@��Ӻl�ZNL�j�z"y��&��;eۮ^Q�v��'�K�"b)u��zKW��*�QN�2w���,P%&���l �p�C�Q
 t�Q�-0Ļ��/{.���>N0�P���ۤC�K�=̦�h`܋FjR�����%��닡s�����MÈ$A��F����r�¹٢]�]%�GL.x)�Y�pe#�l��4��ɋॉف3ʳ^y��Y`�^~�U )R�����ҌT9�hA�)�|�5[A�(.`��tܙ�W�x�V�(�&�A����M��I��
3�
�8	֡bl�V3�ZJ�հ6�T��<)�]oH��m����$�U=�UI�k�-��T㒵+?c%��R�!��Z1U�rxHj ��i���K�$V�c-�o���z6��A�T��c�]��e"�u��z)���?G>7��fÍ=�¬h�="��w0g1?��|E���}�MW�̡�t�Ə��̖Q���ұ�`�E�������٫`��LUMQ��Tz����|�Ô2}�V�-%
����6���"�ⵋɸ�Vj�ަnbj�ڕ3b�ەK�uHC�z�����l�a����m#,�q\�fJ��� HFPEF�]މ4r����������u='�12�����F�A�602*��)��b���s�d��a���q�pez|��92@򍶹��CK�<yr�R&7.Q� ��o1=��c�=�f�iAv��%4̵�{
��\Y�zPp�煽K�;۪��O�����>��dB���C\$���l�]/�p٪�=����]ݲ�H ��wA N��@�ԅ�����l�L1T{s��6L�U(ϒ�u����rb)D�+�x��L�HJt�nX��`Z�M^�w�Ŗ
�g ��i��1���*1�M����J����ؚ>��=JO�-c�\��i��� ]��K���S��j���vr��� wjl<*a� �88��:d�T܂yoj���2	�$xyݦ�6w�hM�+���v�%��C�Z��\�/�T�j�E0un]�?��<��yk0�ʴ��	4�!?9�Qql�K��Cf��{U&*P�xF�Ɩ�S�_�����������CB�,%5��������\��j���q�X\�?�8XUǥϨ�Ǜ��BGf�/9�m��5^4��'��@��O8���ܛ�WͲz����6R�4�m����;��2c��E��y��v�ƴ��^;Y��!D�ۦ��j
�ƚ��T��*�	A���3�e��I�|?�����ζ��2)9�3��z��뻃S��g���o?�H�i�����ȥ@	�g{���܅�L�YЧ���V�w�r����)B��Z�葞�řN�E}�k��=0#t�粶�)8���i����ˋ4������ݮ��ʆ!�([C�T�����5�o}��Nf��܌9Voe��LG����V�h`�+y���>�`h���C�S,l-���T}�@9-.T���\`G<��\O� k8��0-�4?�`��	_F�X�ׯ ho�)u�5��*>�X��[��
�5]]|Xs�\zv`L�<�⻣�`�_�0V����.���O�C��?[þZ<�C�4��s��iw�F����K<h�3���H���ڣ-��yC�i����^�;q�t�h���ʋ�$t(��%�����	D�N�Z�0L>�E+�#�|����rzCC0�Y��*��6����뮁`�X&uTCiAS�VI1��W���UȰK��=|WL�oo���k�X�6GV�+��uOd�)��JJ�s=�g�2?�b�%u�z*N���s]���1L��g����������h��.K�=�(U�<��SբBL��s����k�!^���?��*��0�2�]E
������@�SY����n�*�SҺ���Z�A��:�|֋y�����J�t��	E~\�]OZJ�y��f���)Arq�`��rl�
�x��8	z��t�9��~
t�
�v�n�w ��'r��8u�8_�퀷��}з�6V�S��c����8������\�6~��N$S˾J0�l��z�{ ��_9���L��������U0��.�U�ӷ8���㵱`�[5&�}�������m�K��(>}�4z�Ķ��:���91�6���΋)�����
���Q$4(T�Qp�����D�g��l �^�E�p��g;����{3~�0�Nu�������O�dY9�E�*�w��b���2��bTm����_�,�찞d��zr��`��~&��׀���!���I�>��W�A��Io
�j�ǀ���J�ް�;zē0����A;;徝���M�x#:lk�zv���7�O*��X]Ki >. UU��\�<��jz���U��H�,���rV$��*�#^�s��Q'��*]W�@��������C6i�L�u�J��H%'��;��ir�xeq��ҿ �mό�֔Y%����� �5kz)ԑ��B{��g'�8��IX�p� �:���r�8nO��.�JM��iǞ�%����{��{���� �sװ�w�Pypd�|���f����<��W
ڜ��'�k�fx����MF����	o��K0������}�n���'���4\�tx��+�<w,�<�m*F3q	��v����������M ��%^������x��׻cP�M�:%��ǒ�K�]�T$ۈ�EE�8��	Н�����	j* � .�pu��+�5��e��!Ø����B�F{-۔��=�8��գڎ*�f`��^$	�	ٲ7���jR�H9z��Dɉ�k��0	3���
��U9�y���'���������v�c�1���cfQX��f+c^�gKy�� �Y&CO��u�W7�M�X�������|)}+�їڋM3[N�aw���#J�φ8X$ȓ��w#�{\S�#QDˤ����M�AT�߀�W�KB[�{��>�v(D�o|�����%5M'�������XBq- ���md�0}��Ā������U���(�wV�p�$�$-C.�_F����E��<t�ky�@����rS^c��J[u+���������?��Z]^E���7{���Q�u�ڪ���dc1�E�x���t*x����+�B7��k�� ^NI8�#U�����%rYȤ�7�4%�[��xN��G,�W���h���؀�A I��ɱ�UKS���������H�+|�Qֲ�H���o�e��������3�Mv�Y�z�����Y:P�ZŇX��x',�Ϝ�k3j�[�"A��:Q!�C ���WєQ,"~Qzw����/h?�)ĥ;r=�ͻj��+��������5E��grSq���8������J�<�4ľ�AO���]�~K�E����C�
���wV1L��GMսe��iи������2�>���J�)I� gr��DHM���Ǯ�oT[Do9�X#YUj��'���w��E|����w#p�>i���]����
��{���P�� �˲�^�̪H4�0��N&cԫǎ5i��_׀�� AO���ݰ�,��2��;(6��iPޜ��|���嵏A�NX�=uͥ�����1�@��g��������>�z�V�I�X��Ϸ���"m�/��B*�X�E�/ � U���(�2p*�x����:9+��f��2Z�t������"�W���Cn\y�BT�*s��j\k���Q~Ú�{���0/A��ŏE:��?s��u�Q0xYN

5���,(�7�w0���T�C�M�xUxoI�O�ލt��Öa>S w(7�����z [�س����X SA N=�����-��R�N!�&zX���i	Ύ�]�D����m��� ��&ܝ�.��@ݢp.�@�*x����5�AG�r��=���6����!�[��|����y:����F$�#�G�՛��!�����h��f}s��pؐk�G=c��s,�ݒ��B�\�Aey&��0��O��Xz�7-y��mH�3�I����=r���EYt/T��y�'�#�~�b�I̅s�	���W_k�z�T؝Kl"fV���S-1i	%���)D�Я+��:wfԱ��@�p<k��Գ� `1�Y�����/���	0�4_0N�6��;��@�n��>����d��ž L��s ��|�`a���T�)�E��y�S*5�� ްL:��x'"�u:��D����s?y�,��"��C��{�����@6X��\�����Ds�LA�
����w��o"*ͰϮ�jt�lH�υ'o��� OQ3��I�����>t�Ɓ��Y�o?�_6����d�Rh6��XC�F2gT3��U�A���jߩb�a��w��0gtC��j����i�������xb�z ���\ڲ]u4��U��p���YǎQOX��|
k('�����.�F�����v�R�tk���Gr ��Y��@02]�|=����D�� &�S?R޺���Be�F|8��;A^Ir�s�$^Ec	w��{h�Q/��U[4�����ff֪���7�6�Yh��#Qh���U��1;��@ӆ��z-�ǫ�N@3�)�������҃��?u^�&t΀Uۼ�f��у�$� ��֨�1\�OS����b�r3@�O�t$���A �����8��G�-J7�"�C�)�T��n!����*�:���V��LƧ!�=P�h��h��â�`F�F��dT-��P����졗����m��|0ÄE§������d8�%J�tG����Ř�P>�&��a���z>>�X�Dp�p_���%b!��vg~,�	��7#��'�D��8%��m!l'���͑
S����햫�`]5�#�-��6�8h��+���Ϡk9'���U�
���gF�L�O�{�y�)\Q�g���!��hN�Zj]+u��d0����Q��h�<�9;�ly;D�L$�!�h��9���LjC�b�:�W�Q���R������/���������X�d��?Y_.Y��v��*�Z#0덽m�
^�b���au���{�8�������QIzr�����^�v��(�-��Γ/���6����$��$�b�W�Ol��=������V��1�]�4ھ�����8�v��i�����L$xw���=�T�C���v�K0}�	��*���������jO�p��� f��#ˀ�Μ�c28�@��q�-���/��6���tA1�&Wijx�a�/���(S�'੩S� tw����|&h���V֯�[]�,�q��ɷJ� T�/�X������[-�I���~n.�8(�꫻��o-��0�B�V�s�>,��Gx��?�<�Z�>ˠ�oiն�ޡY�|��2͎�����6��[G�h��F-�ц�e�V"5��^/ѐ��ƙh��x?��`����}�r�5���K'�Q��v��:�4��7��Ml0�A�jS���8JHIڕ9��j��epM��w�ޓ,�,KOd��&\�23J�b��������� ��L�,1>z6�_=T7��4k: ����D@�"�R����m�������a���X���"�yn��c��t�Y*���Lu%GgalM7�7BATL����~�(��έ��<[u�{=T���3�)󀆇d\�r�Y�:a4`ҋ[ 5*o��I��1�}�us��-�����+����l�i}E.K�4K�<�Q�I�^���p�4���2�p�b���j������f-u���F_���p��%X�j��dpa%Y&>�c�k��ٟ�Q;��]Ǵ:�ܔͼ�h���|;�y�1,��;�Y�����Ⅸ�2kn��4����������XKB��2�V��g��3Y�H���f鶄\!���UA�/��X��U����<�^�#�f���K�*p?�$��c4�ãz�/H�L�����`���I�4�WӃ���<&à���_���Eؑ���_�Z�I6�e��;U��	���rY!�q;E^ʶ�}���iEE/v���H���:����`�� x�
DW"�?��������S��`���+U����
7�iS�.������69Ci�΁���c����I�y��AT���?�-1p{E��Ϧ����⻭�3����� ����R]� %�����C�8=���`D]C�u�I�H{�'�-���!�R�I;Q�?����!���<9gO�	Q?6r ,�b��	n`H;w�����ޜ�_9d�d�|�ܗSO���x���;jfȆ��jei���RD��N�OS��V��sn��%Ϗ����3��n��eZ1�U �R� ��@Z�;j�PIz8��a6��"\2�h�mP���������� �3���ۇ��?;�QH~z���q����(�4����{��%�M��@I}�9�h��~������)��7M=�P��ǒ^��%بv�/=��I^wr�<(�27�w�w�[��І�w��뻲�D�q*Hd����">������~��y������G��i�,2\�h�"����g1�\�4��$]��>���,!�o�6��#$�dgi���-��)?�ӎ��6^�ܰË��?fq�\�+[f�^+ُ�{M����)����<���ޖ:9�|3�%��2ƺ�n�U�E���*:d�x@g����=�����N%*`#��A����g!��?�˷!@�:�h�1d�O+�g������RȓC���s%���xN��'��(�	r=/_�=E����K9�I�1�#]/��!�H??������v������_�k��]������yop��'�!5���8ã%����kǓ�8�k��#O�[f�Nه^�����x3\��ji���V�B�:��+�C���*!9(��
Ϟ�˱I%;1�!LK�{.ӌ.�o��_Yp��f�QaK����!R$.�Y�1,X9���dUT���:h:Bˍ��e�t
Q9	�3Eq�-eQ�#c�V?�Q� 4�MX����Y��>�S�=�^�f�b�9���L!^O;S�GhkP9+��j}����1\1U�=���Ҕ�a<n/Ts���%�c�zT�YW7D���/�� 29���Ic�`f:kβP�nD?q}���n%��Ҵ}��C:��vj(����������I���/���%&����[�%�(�in~C�\%U�+t\���Bi��%�ˁw!w.͈+�Mh�a����t�l��Ya�V�v*��M�
��)/ق ���#�p��T+�޾�9A�����~�9���DU�~�=r9n ���z󍏛�r����5�ŵ(�����g����S�X���.�"��t��]ZX�I��U���;4�S��-{���-�7���ֱr�H��oO�]�?�$Dt ���{�#q�D�����O�����! N7�I�=�D����é�<&H�뼴����{����N����Ѧ���jn��hQljk5�b�R�#��o�J$�F�6�g�+vq|g������!��-I�9��y{�6��OƔ���r_�})jK4dy(��TD��_�	rr=�RM����~}��G�Q�:��G��2lo����|9`��xS��b�`��л�?�A��������9jj|��$B+4���sO�6�L��� 9��Q刘�B�. R�Y0HPyJ���]��2��t��dV����/L�}�(j�T������"v2����:�@��B7Tu
5��r������V�|���H�.��S��	��5��c��.m�^��m~���&�`�+?i���nT]V���Hj�B(/A{���i�-�t��'2t��p�r��)*�-ꅜ�4�<'��L���x6��\x�"!}VP,��x�(.�j��o0��aԸA�)������?9��`�U*���ɕS�6l ]Y��h�V���?DVV�;4��D�C˶����R�{	'2�P�!�����{��A'�jG�b��=�f��;Þ182���R�����ї���UP�!���/=v~�3p�5~\���$:'�����w�sUP`�ؽaZs�>?=�{�_���� dM�[s�����d�9��v�E��=T]�i�[C��[`�Wv �J��^�.k��yt=4��Fy�>�ē%�.��1�@S�67kSӉ.#��`�Rt�a�/��Y�R�v���pC�Ƶ�JvX��9�LWp���\�
[y����d܏+�E�Iy����EOq���o}ڵ�$g�;�Zc�pi-�w�u�Ⱥ`��t0�E�8d��/�[���?`=�ϯ���]�il'���N��CG8�]�`�Ri L��[h������]D'^w��z����2t��l���ƥ�Ʋ��[̥q�`��>�)�$fk���Z(���z�M3�|�f�|���I$~��ϳC=w$>�;kC�c_��g���l�///��UNZʋ�ڡY��_��/*ޔJצ���&���s��.��dQ}�~#����KG��PC/Y��G�w�iRq��L(�����Q;�:��@+Ae!�M�2�cL.��0�s���O��(eDuL�nnC�ˊ�\'���R�t}sh���<Q�@�X����[�H�6/��L��u���R���'�6�UT�e�Ri�P2���rv�"����_����qLW�,��џ�t��u���qo,�-�	�C�L����+g���+����]1�]3tJv�'�"j����ud`��)� �(RT�A��l�~�] ���]ͯ�M(6���_ڀ�9;�ƥ�b8���'?� �������G�BY}��Ӭ�������)w��e��syu�y��s:���ֻ-��0+
=�}��J����%��,��R\����S��Ʒ� �+���o����r�<�����\ߗe��ȵͧQ� ��&tg��k�<��p��y���������]�܆�F��pe`��Ƶ�>��#Vwq�~G�g��!<sw�.�c��֝t�7�
p:/6�5p�~��Ս���<
?Բ2�~�##/��B�_�K�>yq��ɇ�@�q5O�|�%���f��=�Ւ��É0�s`�g�hJt@�}��(*������j޲㉘�4ҐX�3�=Da�Ӂ�H:K�gX3��&mB�qe�i����%��|��	y/nsd��ia�Ɛ�)��lj�Y��7�k��|��*�O=2f�4w�c��B�J�� ���-�CMs��±\���\���s�l3^���c�XWc�7An�|0n+�>�(��^�4�Bz{l�7��Y��PJ�q$����mB���0%�22��K��I�I��3Z�Vp��<.q�	��ch����u������l�r�u����e�bv8E%�;�U*�Z+*��xAK)!'������	��9ot� �ƒ_��~~h��N��Go%���04j�`�<Xx4������Y?����a'�`v�����A��pLl-��Z�F"���1�(�*&�?�a�p7:���)�y���#i���M��/��Dj,Q�A��`��9��'Ѐ�.W�&mO���5s�I��3Y��5+T�Z^��ބ�O��(��n
V��HC�dC�!e�S���zF��D�C���f��c��VsT�7;UH`u�~��E�g���7~S3\QD'R�9:�
�/��e�D���l"��W�v6��n����xU�g�Nm1�	ߚ�-��؜��^���y�m�����Б��?Y2�'�%y?�]$ &#nF���'���%B1GAbz`I�*�{�A�M|�u{W6��c��~ 6�G�w߾�u����M/U�u��S��:��(ʺk��?���~�b�m�B�}s0<D��ΰ"��USi�b6�r�3{7r�%M�,~�ڻ�^H~��47��01wX�'�g����+P��;�S���͂#��]���q�E>P}�u$X�7B�]�&`�
��i��s��v���;Z�����
)�ډR�Ԑ<��2�"���[7�GyH@�B�A�`�0�E߭Y��r ���w���	�15��2#��k��%R0�B	=��̝�,�b��o�[M���4{#6_w;QFT\D:�p�M��$�0�Ș�d3:�(cL�*�1��� ��Iq)��YS&O�:��@9x�
�luoRH��1���b�>���7�ם�{��j��_��˩��J��x�(1-��'r���Fª���w��!C̱ʑ�о�;���L�v�:= �t��-^�0����wk���'����bH|��c�:�ha���
k[�?��N�Ɨ`�8�p�éT�b�u�^�K�}�|`�%CV|��(���� �C����U�죂�/r��cq��}��L�)�Q�5/���Q�~t½ ��.ߞ�ЈΓ��4���͏��)��;�bwɡ�����=mbQ|{h�Z30͸��;긘�Bpc>�ֻ�f�GLs�,���ǝ��M#jl�4M��Fk��x�;�>�Ɠ�Y
K��%����f��LId���uU&�t �����xd�` G]+/����m�=0�u���x���V�n����,���$[����0�̓�s��jL�� q���D�~�I��*A�PE�G��&�a.SXɫ��C(���W�,�m�	���w�"� �a�Ir�;u���|��u�3:k�{�;���P�w�M�k��v��� =�H�}e�ˍ�C��	�|�WC��q}�@�UF#���7��"��U�S�޵_2�iv�7m�4��U��:��bf����n�D�"P`Y���el�5[���'�c8�[}h���	<��>�e&m�8���-��1��P�<!��x+V�����?�j�(3'��	�W�da�"Ӎ�w���x�pIm���*a�e I2`1c���C��h�].X��|d8գ}��Ak�ڙ�GƸ)��k�
�үJZ�f�>�č3A7��c�ŉ,ƌn��H�,y�ǋ��/��Bb����+���Oͩk��<"u�bU�%(�O�24��G�-��3����z�ǅB���oD��T�c9}�#J/Ť��Š�*��O�����&
 ��;A�@܌�}-Y�!sO��M�?�l�pja�p�H�����:â2F&��x�5�o�$��}U�A��&�	=�B*�5aG����ɰR�$H�o�fd�EH�2P)�O߼݂hk�ڂ[))� 1`�'
t~^�4.����Vu�fE/���A������!���@w�7�<�x�R�D��;˙G�r���X���7O��6��dvm�9��k�V� Q/I"�?8�J4b�eR���!�8?칄�;��L�5��;2�R���&�T)���Z�m��yt|��eJ�j
,� �/p�/k��w�N.���u��0�LaQ9�Y�p�gӶ�n��5��G�%iy�{�*��G�]c�_�LA��"ʔ��gF�M���N��:RT���~·�g�K.L��:�"٤���TX�İ  [�+�����o��"}Q�����n^&�=Y��n�$��g�����y?��UCӝ>��'�d��Ò���1�l�w��<���6+/��E��J/Gƌ�0�V,�w���q��g�]�Vh,�|Շ>NV|�7H��*��B:�58򨥼t���w�$0l ��V�
K�&)Q/�?��.�,���
���v}����tr8�/q��)>Zm�֕Nj��>�U�OɃ=��H����TwʴG�R��%E����T�ا�A&�����Z���ޘ�(�c'Y��eל��j^R��F���m����	��-Ұk2RG굟)$�8�\�����t�\g�5��6�҉4~C�)Jp��o�\�1��s����Ҧ��f�@�}��#���,៺1�����x�b�u�a�2������UL�;�f]���]G�I�Ӝ��ѓ�/8��������8��{a\"��,�D�E���e>����a�`ƫ��i&���զ��D�Ȉ�G7n��;�ǻw�\�������k?"�x�3�nq�7�,�X�(�x��m�^�@]O�-����ͥ]��R���J�!��ؐ���>>�2�>� �0��ǥ�eM]�M��i�T�I?>�D���-��s��#xʅv��2�e��%�)l�ôu5F�+�,����k �h��?�����fI�K��+9e��@��]�Ij���M��W�>�y�z�*������Cp�H�~���p�F�׫�w�ɍ����15:Qzr]@lީ�J��%hp�?\���Z����DB����|�R�!�M�1�T!+�<����6��X�͵AlCIM�Z�*�[o"���|f�E_��䶽��g�V���_���Q$�;�p���K�����y�[�������s�G,$�@l~�S��U��2x݁-�hܻ�ty֐�/����Q%<�d��Զ:?7���@�4R�;��:�.^-D}.�*��*����}��w��A����С��6P`1���Z���9Ri%&��L�,�n��}����{%��2��'��=@f��b���0�*��=�z�!��$,�C��kg#���+�L���>�⮈8l��Ó�]f�@�`vzMzH���ݹ�R?�nei���������Z����EdW��#��!�(-
$f�"��*3VU�J$H�m�!�h�3l]��Eɚ�����X�H#H�b�}]��i�2r���n���Z�D[��RZ<�{jh�+͟�^��O�";�ePs�l���Y�d �8M���Ff��Ĳ�B$�䜌{��IF9拙�^�Ƞ�{��HܱN�+� ��l_�Cj8	�`c�`��t&jH�p���~Q~/��|�Ҧ!��=�H�#(����t�y�b;��mc33W�p���tF�HS@�S�
�z���lL	,TkԷnG����'�PT]T����_���~�����l�lb�W����Ð��[��v��f��VV
���R���4�Iu.��ʹ����4�e��L��G�I���$E��vD�O�c8%&����(Ø:��u)z����r����-{Ԩl�d�%!�ݱ*���HNK}; ���7-e*�ࣇ-���>mXe01|�IMJ[C����~%�@��>��C]��eѐ���o��
��'e�8�0q���k*��^=�	�T@7���Ig��訪XV�
��}0� k[X�i��6|�F&���8e���ݺ�y������/�Pq�I�.'�WK����
0�˦=�/,���"IR��.�ǟ�W�*!�-�McK���Og*Ԃ�ڀMl��uB$@A6`�}������W�.%���?��9 �n ꔕkc�l�v�`U��]u���-����N0 �!�Y"��P�ѱ�ph�K6���P1���i7��)��յ��mMo�է��Neڷ�R�St�hh"1�Q1�O�M%�0O�r�g�K���~s8�5�J-tQ3�8��W51:��L�6eE?:�>'�He���^�
�� k�@z��3��i
t�p�\�Qe�5�P��[��Ҁ%�Bj%�	��V�⺩n�
�W�q
��Ѷ�F~��EsU-��b�b��>b��`��|���չ���Ŀ�jM�L���O�&�7֐��6ؖ�7<��Õdp5��6*&���K�XE�^i����"�m.i�{�q��U��?��5D[�⾋yr ���nro��,��G�~�po�M����Gf4���6"�xNR��ju�\k���1��h��?���ꖟ�����I��P��1��&��n�=���5� ]���W?>Uw��%G���mS&*;��+�C��7I���~�#������<݆�� U�p��9�%����	�#!�/}���}}	���9�6S��>��(��bmž�J�X��:��K�@j��kk"�zq�. �4�}�����7�yw�7�rb;�1P��H�&r��&��¼;�+���.�Eq��HE@% �����6����:O��T���$5�}r���z:�>�6�H�j>�|sٺ�gΛe���?�Y��i����	&��"��:�p�r|.�M����wz9�k����Kʱ��U�z��Ɂ?����*��֗.����ZQ_j�:˵38���8�Y����Nض*X0�A�n�@@Z��ȵ(�����.�"�$OQ:�	O�]+�*���{ [Jې�0hy��V�
�,5ѥ2����K�R���l��� ��ƛb1N�����w���c}õ*r1$Drw�� D~RX��n�1C� ����Xi�蕕#����I�"�[y�exPτ�dܩ9�7MJ�/1�ƭGV�{�
E�������K��o������X7C5�d3�׳\_9���쪀hh���za�L��^�	�	KUY}8�,���M(խW�GȲ��X �5�t$�h7��p��r莊��L����q4�`������Z*��T�;u�V4�xFR�U9��V��_�� ȳ���
ޭ_�;��N�3���=�`�G��r���60)$�w��2��w���v=��v5k�UV��g���x�T�Uyw�YT�n�`�(x�s�{��N�,	�$Λ�%���D�@Z����`�Ak�bh����=�������4w&=$I&��u�0OAˈZy%cXz��B��fNv~�#1�QN�(H�F0�3���9��Ķ��?w1�N:{�8F��pu��z��q��sU�b%�z��k��V���xݸo���hU�JR�B�QS?b�_j7���>���Z���W �q�ð���N�Ds�+`�{I;U��� �(�3�BB��ۼ���I���T���!
<��J`��A����B�� {b�hT�>��#s��",*�v^����x���iu��>K�F���vqf�9]:��J�6�~t�
��ۈ����Q��a�e�<�A�sI(�H���zPl^fp��t ��Ʀ�	!���5�#w�P��p�����&�A;�	��`"]�����7���p1�շ��B�V�W �I]4�lǾk��R��t��3x�p�o4��=1m���;�s�^ŭI�a�I44���l�����i��o�������_q>ʮk<����ڙ2��qf�L6D�ugXAFk��5�]�2����
��I���r�}k�w|���H����6_7�
4�Ϲ ��w~:^���4��.�/�	v=�|<w�c�������ߵ���D=ێ���9?f��O�@���i��
�;saT6γ�\�`c�Ǟ�ݳk��BhȬ�ϱ�T�(ʀ��V�0 �C՜���7�A,u��[�fT���U �L)�`4;����Dx�� ��Ѿ�b���-�unQ�^CգI�JA�jܑ/��L��A�?$1� $Đ>������]���#ODR�O(.:KQ2
�D�d.e���J��4����M��_��� �܅�U
�)W$���E1��~^n�Wm��:7U(�;X,��m/k�G���Ќq���ɗ��k���M���ƈ����3��d��5�7^G�I ���n�9Zz��n�*d@�nVρ�O��T��D����i�rZ��U��-�_�%�+ƌ����y�xd�t�l������..~N�����2�cS���GDz��}=��l��X;d��7��B8�>���?O�g���f�B<��Ý���r7L���(`r�����A&r��Q|M�"�M�n[X"���sê�G�b��ش��������=j�&�)�g#�Ľ����� ��5�
pSbk�ɟx�\��#��8�Y�n3�M7�x�%�%�J����W�_����u�pdϻ�/�R\���ulA(*�����!�r�6d�_%��g��"������n��Y���r+����"pV��8���"�HS}�����'�gP'/�9\̮�N��0��ӯ���
�@�{�rۻ��(@��Te%4��d3��Pt�qML|	�k�0�U	7$�q9n��]��*��\�[��bF�."!32�H��������xv����āW�4nʃ�Ev�lNX���/$����vhu��\Q�������c�Rc��UQ۰<�}�<M*�U��Cj��YՂL�	[�����0R�## �-��*��
	o� ����)�k`�`&[�*�Rf�c�%K����X4�ܛކ�O�����#*����M��{���ѹ��OE��AZT&�y
���t�T��=9	�c��d�;ue9͊=w���S�N�:��݋-�q�^�@:9�~�	��k\9�[����k�..�x���w3An���h�>͂� �aGr�?B������fE���ϐ���Ҳ ���]�"��e��0^�R��y���ӫ��ˤY��h�R��]`���A����㢯̩�rr�g�;���m����0��>c��7Dg����x�7ؼ�k��x�VU㸫qT,���{9ټ�n�%^�/6B��w8���'ֿ�J��7�r!@�$��eI1�$�OkVpXVò�m��*���Շ�R?��ȫ��x��>��9�Z�A� �a����=�ڬ�����}�ڳlY���b�L�,ƃj�ҝD�>������Tt��8�W�x$�'�P�wh�_�~UP����*B'�� �w����]���P������񈸏���Ӿ��(�M��9Rf�;���u`����G�X�7=:��������_�m����I�%שY�|� �ɣ��nwg�]��W��xb�-hA|�������w[�-�2	D+��`HL8E���*{�רz�.#�|b���t�e�46�>,<G"u0� Mz�IKB;�u��f	��8x�g�a��v���y��
�B��TNW�d%���>�(�T�́��;�-�D��6;�OC��� +�20!�zc\�Zjv�}����/9F�������h��-\�K&c�*�<�����]�7Z�/���`�Dؓ���5��&x��a���]c�1n����9�Nuv^�\�V���Y]�p��6���y��Q���(��H��|I�����2Z����6��<��������v!���MΪ*Nv�x�ƴx�F����a�nI�_����&�ޤ2΃���i�k�?
�qx���o�&*t�[J"*��n�e��Z,�g����F*��Y�8e���qo!�Y�{�8BM��ǖ|K�s����)!JB�5���������s�%�f�2�4D��j[�vq^n���u��U�lo%�.ki�/H��RnY� �;�L��#�2�T{操@ښɠ ��nǕ-wЯ.����� �{-g���n�X��;6�U�Q�;1Ͻ"3��ܿ���2��@y� e��\P�g�;�ؤ��yCI)��q&�TTuj���J����:��I��!��R���:���	��֤g:	u�UM�l=z�=4�ޏ�ѱ����%Ch4�"A M�?@OZ�p�Ħa����!�G��e&�c}���\��˥;Xj	���9��F^�3$#��*]m�=�^yd»�4��_lz�5x��[?��;��==��l�>`��˥��p*�IH^�Rr����b�6�ϻ?I T��Mo��WV] �}��"Lfz��W¬ )��ֹ}�+ "5�O/����M��d��9' mu�Kd]EO�>���,|�_g�~��a��e�>X�޽����V�Ϗ������
�ڝ�,��0�`�ڣ��%����Z5{~�Ł��s���?�U^S�n(�6��$G�&�/�{ �	4�f��@S�,`%?�Y�M$^�.1�gm�~Q���_K�V�iF�����9��F/�S�͔�����l�0�+^W��������o���O��+e�%g�7��0����s S�Ǵ��);�����=n�ڿ)���~�y��.��w��y����k�������a�a~�oz�a��5���"�(�tk;�����I�bvz��2jb���f�v�(��RJa��du���0xf��b��貃�j̾�׼��׮%!Y��,a��|��P�[���i�U��H����y*�#��P������z��_n9�KlTP�e��#T��o-�,/һd��@��Q)��jhP����8V$sH&kK�^Y7��//��zƛ34
,A��e/�C�n4�$R{���z�i�B!Ё(T�	8e�������A�~2	�柦�=J�}�Gg�[�҈g�B3��,(i�&���)0Rz��9Kw��A��y5P!�%�=^�w�여��*c`�5X��ee���k�\ʿ;�.00�톽�j��'e.gN����M�E�����Q�s5{����6QeJ�NW� �K���2���� /�\�b"Jf73E����|���\�*UZā��Le�xz�f�v���h
��|�u  �vS����Jƚ,	�X؀�]�w�C[��nMh";,|$CCRO�O���7����Cֵ���=���� �:�c'��z��O{�c[�a��^a`OP_SNa��'���m�p���~.׺d����j�t?P9�U��C	sʰ̓��� ��7�F����X��5(βx��"䮍�� ��"	��`U����Y��o�'8poӜ�ԐH������0��n��H�:��W?�5��A�:��H<���ٮ����Uu�k6�?�m���1@̇�ΰ!�M�ں�]�1�#p+��aOQ��ᙄ�����i���REb�AC�4����DN�	8f���[S ?�EJd��*�pڴ�<w;&���w'%r$+4�R�*�����? �>R�m�u�����0�I"�Y��l�(]+bQ����}EA7e�,<%Gj
����>�.��S�\�a��U'ow���Y�<}���yS���3���Ѯ�6Q�.���t�gi���V:�ӫ�<������iiђ���2����Y�ȹY��Uu�$�v��\+�k��B�y��9�?Iݦ���<%��} r��l���m*�^A}��!�\]��ۗ�`�a?�;}�.S�/2�C(�YB�t��;�C��V��7�"He���8��n%��C�Q�\���Ǡ���~��+�z����Ft2ː��w�uy�T*�[����P8=����^�H�Z�%��8����$m;�ſ\"�U�5"���o�#��HX�;�N�V�]h���JIM>�$��+�__��Y</0������V�w�� ]���@D�%Ho$��p�V}Ǿ�6�	k����a�dp���Χ�*����H��s�9�<K�v�>�)�,V�Q,�iV�wF�%�6�wq&����
Z��"�W�a)��N5�zO8~w��S�����X�!�A�d��v�P��_���]R�fGY���|��oU a`�B3'	��Rtd|����l
���������]�z��}�ǉ��,=ֻ�Fb'�euv�`�C�n�M�n�l;�*�ԎD��<K�2�F�F���L}�#�f�b�old���Z$����	��4@ 5��$�z�Z��\�׻ϗ��x��6���]�Z^+C@�d��}���lo��Wf�N4x���-$OF<S��Q{�N��G����h���_m��!�#�P�(���1�%���sL~W@W�7>�Z�b�[���b�ƞi\c6]GN�;l 5O?�P.�����F�I�u��6�,�1M�������WW��X���q��ǳ�9(aSN�b��Qm�	߀��mю��u�|�\I�o�%������g1�|�sK��|2�s��i�x��'Du��O=8V�ۯ�&�'F��yq��q/��(�	n�������
�-z�L���)�d�&1���*ɗ?�>^u���E�|~�ڨb��ƛ������i��3?��_��>�U�5ҕ+�0���#NϮ9a��G��i�o�4Zy��
O��4������-\��ƿ�����Z$M4.O�����R��{x�f����Eڦ�0�m��)d�i&��Jwp�m��~0r|��n�H"�L���s�h䶡t@�>"���b
���ڕh�����#A�8,
0�5KI�_��w8��E�� ��Գp�k͎��}{��7��Tm�䜎u�nƆ�\�D�� ������D�̡�ܲT���Lx�2yd��Vh`�K���=������)�j�3W�I��&,*܃ �ޟM�#ƨ�D�n\��(vsz�n�k��++>Bn�������<[ѧ9�{�$8�e�c�^0�j��|� n�^r��:L�X�y9�o�&����o�Zْ~��ĉ��008Ǌa������^�3���vp>c�fӬ�W6/Rw�׿��o�X��`J#���@�.e��+��4K�N�ڤ��������D^r�5&m��I��C�k�_�JDd�E_�#�W7>�q4�=�&r��\#�<u�OS�x�a\*f��Y�Fww����j�yf��Lc�ܠ9*�}��o3��>���d�ȉ�o�T2�:X���a���U[V^^Q�8���pa`��U���؀:�+d���ل��R�k�'�������kE�CH��6���;�4ș�O�;Z�"('�L���������,���������|�HȏI�f�ff���uD� ߁2��f����`�jtG��ap鱔�U�wO�ЌB'a�_Q��uVL�i�Fj�X�P3ng-���6��f=���U,[��=!�W�� ������˶�"z�x$�2�8#��Ny�P<�ݓF�jòG�\��U-Gs<ڀ%���#O�������Б�'K~`l�Q²��q���ſ���A�j���.O ��i�W4[�P|�� ӰO�:LHg���2�}���;q�C1���Kkwz1�v���6[eM O:D�z�����5��;j#�?�F�LP�J������΅t�t;z�8�V)'���/JNw���IM��y�X�C+v�Qo�=^�rt��g6!���r˜�ɓ3\D4����,��|��h����זN���hO��N|��} :����F�ނ�m��D��]n��%�i�z���F`�p�>����W�=G���K�X����#6D���0�D�dZ�t���6�1�����Ч�o��I�i����Z�2�.qz�;�R�n?IPI������D�e+�N�j��Kj}5�3�0�=�kQҒ�c|���S�����_О��g�Ҩ�]~���z���r����5�����ڴf;���	�5.e�d�ǀ�J@];����q%�G���hg�T+� ]N!I@r%:އC;�W��D/�gE����_�N��^c��.�@�zsqb��hLV{��x��,��3i3�_�T�~���s�$:Ql��g#-hDJ��O1�C�x͝B���`0/�40�N�T.�#���.`U���S%�H^F�d��8�[)t\D]��⡶�V�e�c�W�nv6��r]~�8�c���o�-��' r�����������,%�$�`��{$+̚���K���,�)ġ����[���N�,vGH�����V�KZ��ȁ��[u(Z͵03�|�M�GL�d���o�˜�7V�.(���b��~��&�KJ�b�U�S3��`-��&Es����G����L��e�p�TY
<�/�h*e�I� �JM�K����7R���n��
�#gI��Dx�v �¡����1L�x<�Q3�ϫ�6pp`$�U��� �z�A/?B�#sz����䱴��y9�P8�/�<q��e����Œ|�൤ɂ�:��v���ȷ���W4d{�VR�Ыzϛܟ��ݤ�WME�"��K�JfU�9����T`<���[]�a�=I
ʢrw���'JK�1�9���j�2��x`2�����g&*JQ�Sj+�:Э����j�9���.s��o�m(�uq�,�&P�BE<N�����;_x�ٷ￞����rB��~@��WQE=c?qQ @,�Öڍ�*cu���ҩ����P�r/�Q��>Ď���?�0/���,8��k ���֬���F�ջ�EV����W�����N��Ҕ�yȾ���4 �)�}�o��ټ��~�՛��笊!�����L`�q���.�n�)��ɤdm�P��a5`�*=��̞�?�FI|�՗g3TL}@����#��88�	Z����(�fP����ڈp���`=�Y�BF�����)�����0�<�f�(bѮůp�N,H��z��B��m���z����8xQ�L�
�����B��Q�����Ȇ��1yu�҅�J�>��s�c���PZ{������P��w_B%��u���`|��}���Q=����F��̦���GI�:�g�e05'\t0���wG]J�
��ͣO�L0Qn�xv��i�#���n|��US�����_|��D?A��1��Y{E>��5T�E-���m�Ѝ0���aj_�[K#����N�b�\���(	�f`�s＊�5�-IX���7����_�Uv����C��2�kէ�,,8�x�'��zT\��]]f���8�2�(�����q����	53��S��e������t��4�S�
��'���|@���V��Z�}��,n�@�y�W���>� ߠ�P�,��`vM������A7XY���`��)d.P�(�7�qwq#��'��^2����쑹]i>]i*-a�27L7�� ��'�0-3d��tL�d3�N3y�E;@���G�[�X���j��@5ш&:b�Djӷ�`��FȔ����ox�R��`�#��$�p��9�v��T�	��!�_=�K[q���D��F�����hg"��F���8��/�"���gz�tƄ!B_b%���V�8(l��&�K�;���7�3�ODn�x5=74l��@�8 a5�vZL#�����L���e,���-��^���[ڃՃsx5`����å^�mB�D�S��$Rs!sB$�!Z`�a`��� �� �x�m����t_�_X~� �L���C�;Y�D���c#���v��3w���.��w�u��2g���:�%2 qXT:��6U�O�����n'u��NH8�Aj⡢Qp_R;����v����V�{K���|��;������`fZ���	xL32���0�"�	�R�������
M(�O~�70�
��Z�B�k��?{y	Mq��b��OPl�H��]L�w2�����;��w*��$�C�H�Q,:�|��2�e�@�q��O���k��������]S��9�I��E[�W�,�Ҥ�fxȂ��t$"p��{T�|��MO���?9����2^��Y���w�7t�U��l�q��փc6��s��q{������:���5��?�]�&�)�'R}.Htg t�\(����acAݪ]�W���`"q�|�r�$��)��qՑ���8�u^~M/'1t5�Ѡ�u�D�*��m�t�ɝ.�=�D�q����?+��K���O�����B
�5�&���
��ma1)4CQ����J\�Q"� B��ڠ�=f$�o�Þ��%����f�BR����Ğ���:h���=!�I �����ʜǅ���	�ݸ�z(�}��Kk1�o���'��P
�� ��#�C�sQM����,(�4}L�V|�������4I�5+�����B���א�1��f�f�T�����}��@�#J�I7��/�`��A��
��� ~  ��h���(%�u"�]�W)6M�Q~ +hPP�v*����8�sβTB�@A�(zl��՝R�Y8c5M6��e�$;�r��
�B�ѕh�@���D��1`�wO���n���"�moW��(�:�q������&s��18�܋~f�?�$%��Z�l����mZJ�������1`��oV�'�M�8(e[��a0U�Wh#pXգPf��O����F�^Q�X�tڙ᭼��+�'��7� $��މ�no��Z��3R`ᡖk� ��� �nbI>�����Ce�9-4�ʤ��}����}��n4��� �E��X��?FD���>�<��
m%�_k��`;�D,�����4RO'i�$CA�J����[cl��xr"��m����>�ҊUj3�F.��:���YOR�NC�
��MIP�Hf�lp�C�E+"��4~�O�7=��8�fh:��ç?$ #m�Ƿ�Z�j��j��G�fIۀ�{ݣM'�i~�$\Y���p@^���δӹ(�M���#���P��R�x�ݎ��+�����>N�t��+mu}FI�?��,��0���ò@�vy(9 ;�L�m�Jb��oZ��h(iY�e�AR:��8��~���XS���~@x~�@ωCs�[1ߨ*Vv�y��A�y���"��񫿎�C���,S9�W�1�k[���\�$�b,}��x��ˌ�;P�M�Y,��J���@�
��=�"YIS��G4�Dw�"�ە�>���ͣ�5��V�&�*b�B�!���V��Ԃ��s��x����t{����V0��27�Y��씫Q:6�O{��U������#hA��W>��uk5!�qpǿ'��#��9�o���VX;_֐��F�o���'���j�_+�S�Sᠮ5��{���,~}�[ԉ�A��ܬIv9�pM�"1~���1��s���9��Wg����)7�C�Q��"L��rq2��ʬW��p��W\j�^���!����RT��鮚B��������T��'�)��Ć��3��4�s��:�<?v��"�%��3Q�jB�mj�N(^���4�9v��v����(��z��ؐ\T�1O"���!�{o���Lzj�h��?d�}���[�dY���puw�S�M�B�$뼐p�	��.���w
f꓊ۆ{u���C�ꥎ����bV�:GL�vwp�}8�����Ԯa/��P��۱\0X���$�S�R�p�,�#�J�Z4�$�K���vB��)́Vy������=�7������j@�ݕ���)��g
�˰�J/ŉK�6�U�fn���Ƈ���m't/����"�����r�S0��Sx{��;g��� ��[��f�_���NX}6�y^��~;x��.�؏<,��-�����<D9KcZ�Jw4�n��/�x[̈́��T3~U,ɻ$G9	��ΩLG唂9�{��q�柙�55���Z0�7v���-Z��g&^�	�d4��hu�ab���J���٫=�I6x(�?4�B�-���[d<ˈ�sUG;���*����t�aUg����#Y�.����6�� �B���d� 3o�8x>Z*�����M��&��|�l�|�B-3�2͌�3k|�e���让��p٭B�
�;�Lm��={�񏷒�sUp�yy���*l(��pOkja��� �2vG�D�C���QN��� )�Hk�_j�'W)Hs������j�V�}J�l�@�X��B'I�`�CWI_�^�˧o�a�Ɗ23������N�:�g(q�u�ry�i���o�h���?tU�a0��g�M��gQ�2Ul�x���V�����>;QL`�B��QcIG;��#i�{�@xV4xy�r�W�??ǡOxC]e�,��ѥ���Ux3��룰�&1G��2��í���7�tv_3��@���i�ND�G��gbE�q��#!���48�8����	f�/�fa��jh�GD�������^�
����%`�hm]���vQo���m�f.�ݾ��6���=Iu�``��h��y5��RG���8�֟myK�J��M��b�y��<�8.߆�{�ֽ9�K��l�{L��P�c!�ygE������UN�0U�0g��Эw�$P�م��V����Ź��Q
�!��42�
u��X�i�	}���arv�C�c꣤�JU|��-ẋ�5�%�Zw�T��x��	�ˏL{��H�cy��$^v�D�ɃF\����z��eH%���,(ٓ�aU �ǥ0�N������jg�
���Ls��%�<V�㑸�|߶��8ÕJ^��$ ~)���b�n���c9��A3��MU�v��y��1ΛE	��i�[�$]��{�����Iw�T��q�����|����q)��>%�I�:W3����hۆ�+�1�y�Kw�k�t���0|��j���_��G/\�cH��i?=��j4Vno��u�����p�^�s���!4/���
P��d�@g���G��;9�CA%�� ���ssm�����X5����SS�)�*���I�+����� �);�δ�
�izP�'����Tj�������rtl���T]��Tf�B�yA����������^n���u�X�����o-$�d�%��Y�J�5�8��e�g�{�o���Y��ɜw���_H۱��:,(�"^� �Г�5�~�p�|K���VNܫdĝ�;� �.�;����6]�^�X�p-LEK�r3]6�ݴ.e�%�i����.��X�����Ӑ���I��U�lg��@HT��� ���)r�esj�Ҧ�����,a=�p�EX�w[�,�8mܾ�-����!�cl��Ƚ��1����ή���M�'�����N�uB��f��cLz1�����1��gR�3l6�_�=7��zT4bЏ���L>M$OP�c�H�������jF�7f�	���r��0��,x?����.#�o�
KyXN�����1����= ��WK^�!��*YrTte�zd������6q��/��}�N�1D��5��,�G��ة�.�A-��+8��ƶvnR�w����=C�p*1+���n/B �[ˢ�,�<������[.���OUDr�+�qse��V׵�8XH�{nEߙ��W2�{EH��ɥO��ҟ�x�w����P
��K`x�6D�RF�j�~�HaL�+
<p�=h5�Ń�ھ�<��7U�d牆��(�������E�lu��wKD�M�TȆ��=���b����巛}�
���i�$x;������8�l`LX��v�4g�U���' ��<lJ�R+H���P'(�s!6�g��9��x��r
��5l�����T�0�Zu!Qu|O�ýgK��=�`�Su�U����C
0�WA��$��HQ}d�u�_3#_(�HX���RgVc����a3�G����D
Kf�fE^3���gR#�*֭$����m�5O�|�t�D��^�DӇ3u��WuQ�:�}n���25;tI"��]���ܺv�}-R��ڼ+��������ǔ�@��!�@���ϧ��T�`j��jH���Q/a0Q@�	&G��uc:�G��#��������I���%k2�E���a{E]"�x�S��R}A*�$��@wdS�|�X����xLE����U�t|,�%
v�+5�x��I��
�c� L� t�n%Rݎ��D��.z4H5 ��<�i.s+��6Ȋp깧�� �d�u�,d��Sv�[�6>!�1c)��1q�'/.R^�P�N��-{�=h��.a4{ʷ���5�*��f<�LʹOP�YG�2�Eۡ]f��d��� ���PN%)
N?'�*8�q� L�F�I � ?��[�i�Oe�^i�PR�SL-�1���掂h�o�Y�r��N?9�(xAV{��t)�ʜ�:�V���j�S<����EO�E3p��7HNδ(��}�c�9���\�����
��5m.nY/�ם~�q�sr���o���}�W�?UsPk'b���?�.}�@�_&r���\�e�d.U�Z[t�#���%ʊ�x��������PyR��X�CUM�])�a�/=Zj��:9��{
�>�h��y�W�5��k�t_��$B!Ƨl�^�� ٻDD*���&u��XoPw Y�D���Z�ge�����	�G�!�{��
j�М�]*qB�eS��tk���԰_
�P)a��ğ<�J��	�ߞ/���"Ds�}��0BRӃ��]�%����~nf��g�
��N	x�ܡ@'�"��D���H�V3<�F��R	Y�1[OK����_�t)��fE���_��)� Ƨ�vM�kZHn)v�M�l�u(=��SZ�}�>�/N�H����xV;'��6j����D��3yu���h%�h��v�>ױ�I2�/�=�8���O��`��r[�	:^v����g�v<� W�e�F�k��+���v�ǜ�;
����̐y����'%R����C��R8��tj.���-	�� k���.]5e7�^o2k%��d�ſ�6�:�{�Q��,+T@2�$o�i�qSe-5�2Iw�G���`R�[)����N[4)=��w(T�A���DT&��*K������_HR��/1�~J;U�M��3}+f8+���;�� ��p��ؕ)Fbly	,yjvI�$�ߴ2�h2h-���/)�E<� �֌<��`��nC#?O*>��W&P�!P4m=)�A�l6a�?��$��Ca��V&�Pb��_m����:�;HT���H�_};r�x �4�o����ܝOEP6M�Vt�$�0�0�����h?�t�S��a��(�٤G�j�'�y�$�Ъ��y5�9k�U1m���y��(4�*�d�y��a(���}�x ۇ__�a���E��e�qX���8��t{�w/��UВ��*��"�V�w�C�9iuy!\���9�򆋕SFX*�c�t$�h��
O�o�a�n�~ZGw+~D�0㟢Lޱ�߫r(��!㟼|��d��W�M"�u�v)�ړ����˓�y~s���g��&#'����$R��'��F+�<Y���}%43jǶ��Ooꆳ� r[��&�\��_V1�Q�Q��D���"6��C(h|�ɝl}P��V��OTb9�������W��DӕI!��;��/�p���B;��c�
ߴh>��e��'�t4�dɽk�a&z�D����g����b
W���|91q���m0��U�װD�6��#�#aVQ�U�[��5�<OkA���z�����s��TPE��p����u�T�\
����`���Q`Ν�s^��P���.	��,��ޣ7���9�i�h �;�X��u�|��m*v�e`b��׺����3���t�a��d����5���ǧ�k�J~2�-Wni��on��M���|/vevߪ�D2�-���+�&Mڏ�Z�w�Nn�zK �)�0�V|�1`�HF���;�D.Л�T����-�ܤ�ΰ�LZ���F�}��Ѹ�o�kih3��}��_�V���x�����""WB��6*� ']�Yq�s\�ۚt�$`o������V�A�=�u;HM016ELVu�>�m�q�T�B�EB�������}���!�����(�%��6�,S������7��7�q���9���#��;�u����dz ��.��O��t-�F5b�n~ �,�A�Y���?	U E�)�7�~xWz��`���[1]���턘��?�[�#�#@[�MȣH��ɛ@�J��
��zC0Rs�wANK��s�������}�Ҥ�P�@�������������Yn��3�N{PE%B�2Y��O�ͿH��y]ٻ��Co�]"�Rv01.ֲV�ҋ]����V���F�D秗ZЌ�*5l�����)�'�vqM��En�3��:,�n��|����2��ۮ>i�2��P�����5�`ތ|(���*����1v7�>m�B8��U�2vۅ���B�vPraY��Z(13u~@4��)��y��g;�W)�8&�a����p�X	)W��7gd 4&9	�9.Qv�W�r 2ƣ���<�M���K�К���u`���SU�
*�S�1��r�>ȍ��+��0�\-�1%߸Z�Q>��E���Fr,'~�.o��u�V�+�U����0+[ �(�k���_΂����n�8�T@/s�Q�Nh�3 �	6G�Dr��pp-Ǣ{�z�r�!_0|SԁY	�p@	�R�h���E����<��쁐��G���-+�)j]���{��T`��Cc�r����.�ڒ�z�dt��!�2`�!i�61��KFQ�C��JJͣ48�\CHU��xF�Dz7V��Ŏ�D�N�PC���o��+ 5MWwzW5���mڵ�9���>��`\:�!0��$�%՘J�����0�T��$�H(���{�e��������'ˋD��#ҽ���e���0��	���NI�йR̰.�=R�:*Vy���%̜��t*�'��j�OS�;��zm(w0��@?$W��V�6�����V�p���n�K�"@Mɿ��S� ��] \;���@��Nkz\�$zg���<X�/�14� ��(u�ƙl���j���	�.\�0	P\�i0JxWq��D�gߢ����gO��G�S�Xf��9���Ww��45J��9m��}4�^oq)c�T��ϟ��q�,r2�?��4E^�D:�[
��_w���]2}Y'!	���?O�pj�!{��2l�
Z�[� ���lYa���[�S���Ly8�!z5Gd싰�d����v���>!��m�5��Wv&d�)�4J䐹j|���Bq~��K��(�UM�aV�k�o�TFV��.z��Bh�9�.��I �@(��\-�#-B���W2E\���:G�_J
��'��{�z�у��1Sv���s��d�;	>�������0���N;G ��q�4�e�C���/��(GJ3�o|H��Y
P䝉 �bv7=���FΧXt��S+��O��O�gA=!�VԲ�_x��L�<�t��=ϲ���d���c���Xi�/L��#�L.f�C�Adis�|����֭'Vt�/P�n|�kS�tLM��0<��-��{����L���W�$P"�:��]���q�rQ�\^9w(��Y�+��Y��ݚ2P��T#��=\�-˺�~:[����{:_S��ه�֯I����8������6;D��H"����&:���ʳ��|r8~'����t/V�^o�U�	��So�I��E�����r%X�;��6d��&-Qrۃ��0��TT?��3^���Q��ŘBɩ�P"1�G|���o�Fn��x�Mr��@`F��Zޟ���:�9��Ӑ#������B��#|����Z㍀����c��˅5R��<�2A��UJkV�yk�Q"�u��N��lG�)^�lh�.��z��BfH4���A��\�G�����t� [x�S�H�A�����+�#���		�I��[ʻ96!�)�|�5��ܔ\��`%`���QƧ�<�O^�|��!]k�*QaEN�k�4���M���d1��Y��8j� �(�(B)<:�ݳ�Ar�a7`�b���֗�\��t���a�sʦth��a��[��*Q�&@���k�u$��-�&��̯ߏ�4��N9��yh�~��Q�W0#�Z��)BX�!���B;<�<��Gֳ6�A��_�1غ��Y%iD(�6�C��:PR�nxm:B'�R<��ha���� �>^o�
:S�w������ɸ��o�(�bw�f�a�����0\�#$j]��0�H��~�Z�C��b*H���j��'�s��0�Xg�������M��>��CZ��,T+͑�ñ-��&�g�c`r}�oA�Ki_`���H3ڇ����#Cjt��mq)�0���h��0u���7��M
��R;Zd`ͦV/˖F���Ke�oG$窫���F��+SaE	^"B�]R����D�DZGż��� v���g�o�Tx�bip�������2Z�5~X@�:HS�R7�O�P��p���7%~���[�9Q�@��`�d�Z��^/��*0l�rf�*,����nIx�V6	����]%�12C.k�]G��ۋPAo�M��\en5t ɘ��y��Y7�i���2N��?�I��^��pd&��(Kq@���g�0��A=���6s�fq�*�F�-*'�f��!M���5JY���&t�<>�F���(�fs�e=��Qw���;�B�����L�qH�#0L9�SV��
�jg�$#�^$����S��	P�u�l��w��5���������{I����N�m�=/3p��Q�e�]�`䙅|Dcpf�6"/�T[�35�+ܙE��UjTľd^��Q�������D-m'��	�͂��g=�n<�����B�T��OzSz�j���S~��:C��նd��>sW���q��O�>�u2#��bK9���o*f��€j��n�3U�u6���L(�F4L��4��� D	�ђ�K�6b�~V�ƛv~�?:��3�ణ�3e�Rg���(߱
X�i��'�r�@�ܖ%�Y�}յ��G������+����s.�>K!��Ȃ ��q��"=�ޡ?y�*�xV��O�I�����j�,<��#�-5����c	o��;ϵ{p�&a�V��ҫ�˟E�d��:�鴤q�}��a~��
~�Z�^�\4��g��L����Nd��
-�lM.?��y}���8t��J:ǝa�����y����}$�q��;��f�lf"1�`T�dD��M����3��'�B88��Q5IZ��.>����o�oAoIÿ���}{��x.;�˽�a���(w���`[+�x�L�h�DǓ��A��b��P��`��3�ѽ:~(ܵm��<�ҳ�߬hX�F���x���W�!�"9�i��/���(�G�<��N����?h��ݕ'6��O�#_�
9����M��>����������_��l�w'C����'X �tZiL}_�L�u�}�rln����x#OT�/��;���+��t���Fv5�)��� .o�ş=k�~=%�۬�K��E�lsqNm��F�5�q�6��	W�����ѩh���Ds@�-���~���:������ܾ���L��{�E��&fT{d�j�]����(gWh�H������eM���0i�/�
\i�8.��|��eS7&l�\�NuשD���ҧfa���ӂ��0�˃P3�s��aā~O�
����mK1R�L��ޗ��,.&g��,�O� �hs"4
��(�(^�}��-E˘�*�9m����cYs�u��:l93_z����I#��a���<��%�W�zH��yKz��=�������_����K|���z��س��A.�ڕwb����2���m��<��R�3���cDT���AIN �z�I �T؝��;Rn����Rh�������8�-�����r�T �pw�Fy���P���L�g��R���T�%c� �����*����!`���R�󣗰Kn
��g�`it���n����2�x����@x�gBi�KR�\����<�����:7H��W��4�,
��܎+y!�oI��7���<L�*/̡:��+y?b�p m�&u3Z��;��m��M5����$c��D̆�g�7w�#��Υ���v��eL�S�m��N��!��8Hy0��}=�J��U��I�Wb\�Vޡ��i�λ���.dp>э��@V�G'�p�݋ 0�F��E ���Ά��(��[������n���+GU`��<�V�1��
�ϧ�O��u����r�(�A���M�c��Q�D��HsD��� ��.i�m>��<����1���V�:LV��o��$�QL�C;w�����m�\�;�yc�wl������ɬw�Ts�qQy��e.fq� u'K����o��,P6�获A<���[0Y�	�8M#a�J����4�r���Q��?7ؐ�&u����N�;�m��e���s���B.]x�y��nu�uĮ�a������>� *�c��׏��yKz��v�௶�u�
&S4���`BI�]�KY�6?7���1�9�m��m��r��&,�~)\���R@�Y��McX�T�x�U:<�v�IԖ�c�m��Ef-�R�I��7�"F���%z'򉳢C��8�v�|d�?�N<����~�s����Q��d�<�c�zB�Gi�N�\BJ���~˩a'A��-K��Cy���vI'd�$�J'��B��q�X��}*��t���1jW-�l5kh��}gy�3oI���ϫ��Cɬ�O�%*OS�����x�.��@������z���;�$u�̀Ygq��C��A�E�މ����R8�������,i�ݨ���K ��a"��KҠ��ز��=<������Fm��ʬ��!,5���q�d�=�����y��e ��ĵs"ce%�Ίa���Z5 ��>kB;I��=l�IU8�L�hO����w6*2�o:ov��='��P�k�a�ZL��� :�,ws��g"-Ji�$P��#��9��{��eJ�~�W:� I�8�(~u��eq��%X��1�K��9�>	���M�\#K�g1��";�,�{h��a��)������k����|��*6;�C����UAe:�N����y���C�0��ł���Դ}�V֯���a��V���^�R�����YR�ln�:Z�}zn��>�̟�������1���>㸲�6W��4����紇G���(gې�Uv��f��A�메���c��	#�.�<)铞I�-�W�C=�$�asע����B�P��H���%��׃�Eo��@�MU�֋1�W�s�a	F�2�_�����1����i.�P�q��v�\cWjbm���&�w(7�<X�ߦ��,��Q��?|��R������'@�^�$���F�񠊖 e���i�%���U�ø�?�"RQ�}o=|�Cәe����3������� J�v��B\Ŀ�!�9_����zva|�a�Gg�V� �-��nN���r8��9:�H)�j$;��7�pI��d\0#H4�N `#�L��R4�y��+�q�d��� �1
�J4�<C}
7O�kW����&� p�{ypH������K������5�R��e���
5��Q�m����޷�W�h�mg��2U&09.��z֯��Ě��ٺ��D�T�+�̚X�D�r��0
Z���k.�9ZH]�ho87�M���&�ý�*l:���r���]ـ� �:����5�!O�U�VM���Û ���(k����!(�iM�`����$��1����UI���#Ϸ�{����>��}!UB���'z6��d�¼PH�\P��]gj{&˷����j�W!N���d�wK^�����cZ�����kM2�
��}���N�(�E��-�1UC�Oc�
�!ˠ���ϑ�جl�<1��.��ӪL��F�;J5��Y�K��|����QE���,nhg����c�1�IGl�{�-��D�?�e�۲��"�[~2!<*����	xn�&��6�U�oe��Q���n�_̼D��R�
��:h��̧�t*�����"n����jz��^W�RPvt�ä��mI����fAxW��f�bdϋ��vT�Bo� &4�#m� 7�K�u^X�\��e���qp`<H]�|C~�1�8�E9,K���g�#D�}MOw]a��[P�䡠�O"@wU�h�(/�̨��б��!NA���Ĉ��ߖ��	h���$&����T^�8�z'މm`�Sb�wv`�e�E���p�X���Yd�t��� ������$r��:�nW��Z��7�su��LC��%w[�!K&�x-6軂u�sw-�e�Nz�%0i��V�A� ke�54�ɳ� Z��vd�ş�kY,<���L��e�˛/���W˶U�>_�i���������ވ�pƗ�b�v؄�^N��Β~6�[?��/|��tA���muBo�^���gn��%��nD���5����f�t�h��ӕX��#�)�R�Y*�
��4֐�pIY�s��*��Qr�6�_���	N�?��F��I�I�V�
�t�A������C������,�j�6$�D��>t�;�4��D'E�k�m�Α�͛��/�jAk�Yf�1�C8�Ih�A�^o�VWz���um��D��"?�rH��-d\Y�#Hx�^�����
Y�=���yP����*�#�	N�����9-�!M������ۏړnK�P�LP�Yϡ_�D���J:?��A!����m��K�6�{��È\�J!�+�.��T⧖�Q�6l�\\�(�jKEA}�|�!��2����H��!e
�%�h�
��k-�����JY�m�x?���o5Ħ��g}�4y����
�y~�m8o�<��zT����2��PbYcB\@M�haG�����E��O`�&>�0
cJgo4q���q���x�8�qY�;�b~#�I}[�7����y��҅���[���'C��R�� C@|�S(�a��~�)z�ڨ.����/<*��Q'�L�'3b�>�����F_��J�E9��9��ڇ��5��%�)���20O~R9;�#K�t�O��ii��Z��	ѡ�YL^�bW`��7����]����0�����H1�UW�ou����&�&�J���9t�"yn17�����W'�=�,�ro�ii�ES9�UV���W���c!,O�ǽ��-���;HW[B�\�;�`O���N	*�*:��ڳy�K�3��ە���dz볞Pف���ܚ��L>�+f-�l`_&ά��p&�6�����)=�S�A��	w5�_`�M ��7a�C����L�@���VO�i̓�r��U::K��D탬���<�P���i���ռ�����D�yh8^BߘD������Ѐ>!R<�|R��%��X���KbKEú.�_�t��f��eq�3H��#^���2�ƙ�H�X"z���z�%=��2�y���������5M���p�^���*D��!HV�rMsZ{u^�D�I�º�]��$n##�\H~��S����L��Fgr(�p:�ܧG+>��U�6�m��A��v�2��l��2ވ�"�5��	j�IK� 	���5N3 t�5>��ݢ�:�oŒ����q�{$L��=���Tu3�.Z��I�	���v;�x�z �M����11a��P0�N`�C���4	q�����Y�����<�6�Tt���f�E������+��d��`�a�Uaܓr�35�o�����
��)~dR��hdf�t=pb�DZdt���A��v�^�p��AȜ�]O�'n�
r�攸��Sp���XPM{�k\�dQaB�e�2mF9��oـ�Ş�a�5�u���-���k훲@��1ʀ1|^�z��M��]���cؐ%��s��K^�f�|�+B@!����x���Wf���y�>��w"-ss�+��7�<Ƽ�o��e�Dz�WZ�Y(��͎�#�����ѯW��$Y���͞b�4��
���g]���-do�%�M�Niw➳�b���?���l�܅i�Y����Ì�a��vs�:��^�P�|CJ�������������VMd~�L�!�,��"kr�2�qY���x՞��9'�CJa�e�b�`�*{ݰ��}N4�, Y�r�sb4�;��ca֨�U'��T]�~I�L¼/஌��Ԡ��?��0��#ѝ ��q�OܾZ���!���]�ӏ?m ▂�#$2�W���!f�_P^?_ l�!����%�M��K��,'��؆����n�%T��/�b�s��Qmߩ�Ciud��6�z��l���(\,�={��sI!|�U�HӜ�֙}0�����a����qR�}�+|���u	��H�5%G�/Θ�H9���磒?���+j������J����7�O�Re^��aZ< �y�������"�3)>��'rs�����M㽗��l�}6� =�ҜN�hU-���#��f�K���5�i��'��j�V_\��9������-��Òl��;�<6'�	�D��{��9��^?�z�j7w��Ħm���)_5�V�^�Y�ՉJx3UO�������& ��$�[�,c�WjD&�2�vj;�dm�[-�Zy����0��Fe}�蒣���:Z��c�je�ܿ�Coa������e�d,�GP�'���Ε�b���rc�E�>b�~��kd]ɥ���ਃ���aqvW���i����mYh��s��?偶��
����Y�L��&��c6h�0�	eqJ	�]'+�5�蠲f,�4�!v�R�4����>��V�ڋ��oU��Nбvh�=���,E�k`.KTB@)e��D&���
�:��@㹀���j'UcNX�N���L$�3���-��"��du��;�{9���p���w3�=@�-�C���+�y��EЬ�mu#�z�hń�ӟ~7J���f��:=|F!�XqX@9��!�8��a�_E��#:q���x+�L#}��� �/VF뛃���#����� �Q��)
�{y���J�
,k�kݳ��ӓf�bPQ�Č|X�U ��juUV�0��u�p����&Lug��V��j�s\wK�vd	�R�L�9wL�y̎�ғ8�:Y�	�#�b�������jU�,0��	e���|r?oU*���bY��� W]O�w�Z�C���s���8Ӂ���X�"�{�8���uC�!���y���k/,4�\D�?|��l#�,��6 К�Sʀ{���c� OÛ=��Fvþ�sq�7Rkǜ��hb�pH�'ra8&Ĉj�q����Y*�b�=\�ii6p�n���d���ɳ�N�<0ކ�Y�����pq"��eP;ï�S��4""��[���(|7��==��"Rx���>_�Ag����Q�ky��.C��߶��8jDr��5�Hu9���x�y'�7=�>~���ی�J�rd���)��$fF��;�V������4�(�~�a��+1c���c������:�L���1��U+f3����Y�jEH염��t�K��ʼ%�,�nh�\D���D7����p���V���d��{���@i�=��c���x{�C;"	���;�p��~�1����?c�b��Qt�S��H�d�˱�h8�R���u?u%E�-�.WI��9����"M痦81��{"c2e����� ���$Y�B�* %<���?;B�L @1%s\����i��9�^[�[�`�/��/��a��^���k׌�=m�
S^�5#S�G��-��RQ��l���*�;�E���!�~z9ҍ/勸ͭ:&���l��S� 5�֐��$��oi]��D£�6N�@v�vS�KhD;G�I-�v@�5"�9©B�ܭ�<���?���$�Q�6��Ԍ}J�	�@@}�R��( ��XRJ[�R�p��Ta
�h2 U8�,���AX��_B����v5u*N��\�E�6�dL&�M�.|�����DHU��ǈ5�eFi���k���6;���%�^3g�t��lp���A爕��C�D�3��2��&�B:-��L�|s��&�f�x�G�?�#�z���v�)��E1���qU�q�b�mJ7��ƽk��6��1�O�XN��l�,(�p�������.+��
��5��L>B]��!�kZ���.�/K
�H��K�e`97�}�7�� ^_{Ж��jzq��Z�K_�羪h[�ZV�Ŗ��4.0�4C�Py4�0�k "2�0������1OeF/ ڔ�4�.��C��4l�vFK���y���~�^hw�B�h�l�۩��*�D帲{��׃o6N�v��9&�]Yԛ��.L�҂���3�w�w�;b,T��w��!�	��p�GX6���O���� ifu�t4pL B
8ֱ����A���O� ����ffgP�i��RX�w+�C���<V^Ms(�\�~AVj6d"�q (�W��tk�M��<��KMWs���g�S����*��_�?؜���ƞ��}�Ef�([6���n�"�T�1rZ���l'�x\���:��&R|5Th���%(h�ڈ�^d!i�~��I+�n���#I�	'��^o�����Mu3t
~$����75�K�����������X������\_���~�r��$�-��i���ܻ ��S�W�".�+">ߵ<gh���?;�f�xt�;
�$�w:�Hjc�G,�t�Ěx���`y�������&|�4 ��6�X)����Y�#��=b��A20X����+�'���#+��� �����L�����Az�LV��8��8h>��ٍ�5�HԼ����b��y߽UX�;����,@�R0�x�>ts(����U���ɕ���).gZ*�B>���ree��>%�B���f���2eɶ������G<�vG"�H� 	���10�]� �����͵��%쿩��P�h�{��,�� \��!ս"3�9[�Ś�ԍ>/�{`�ʩ�%'�<ծ�(�������i��̊W[GJ~4�K�Xu>o�5砈(�:)�5m�B*�>���o��Y9�
�Z�h��*4����d�Sяj"Lh��o�صG��&mK'���T����H�1��m�GR�D�J���󆇛�+�6����_�i��{�දz<���u5g��=]��PhkJ�I��7�ǀ_7��� %�Z����o�l�b�?s� ��g�]�����3���&�斾R�ѝ�&|ʦ�Drrd��U����.�,��y�/)��Q����6���b�8,��F����bPJ¥��[�BVB���tsTfN'��9{��	���w�F�h���w�X	B���L�[Cj��D��Y8 D��Ău����"kHSluT�~�6��5��b���%;)A���7Yff�5�%U���S��xƜE�A=c�����2Oz� ;�)��dOs��F�S�i¯��A���.�:��[��s�J	�⹎�/�y7o���9}��@�6C�̌�Tx�����K�,h�z
�����l*�]$$��a���uraXtX�����~O��A�ꜥ	������+�f�P��!�@M~�
hgx���������w�H��{�kb��J��P��7q���J�#���-ӡ��D�Z�mqmFD3y��m<Z�	���?����H��{nv�&�wۜl$����2��Qn����[Ol��'�9�k2]��J8J5xN/�SX�)D(2�Sps ���c&��rX`�J���TV��z�}��e���|�˼� ���;��X�;�� &���{��"+W�c��S.%l1����w���Gb��͆��:�Jw� ��~<�
3'����w�'u�3��܎ ����Z�f� ��?�=�&��A����
���Uu�mi&�<�WP.#��F�`�#E-�&/:�,Ѵϧ����><A�v'\<��#�+�0$��}�1J�s5�%_�`f�{6`�8<KB�=T
3�5��ø<l9k:�S$�-�6����F������#��2�瞮3�@�֌3�M:%g�J��{3g��c��~,�����b�uw�({XY ��f=y�z)�Yk6^�)Z�(j̗K�M��;��+�~���Y?�5=�?�$��p���N�u!{bw�����_��ʸ\QBo|����P��#yL;�e���;h1j0k]$�|T:�ԂrFX�3�6����YGX���)�]i=��	��Ѡ��f�SO��NTOz5Eg����J�6���5��spw��K��6U��Dj�FTfR:,g�� �̔�<t ����w/��dW���>a{;�\�9���@탇IeI
�W1x�:�S�oV�����
p�� u��5I7Z�/T�e�W�t��ue�F��a	�W��9��y��M�|M�&-��-�i�)yJ�� 'z����Ps�t,�*�*B��e:Zb%.b�L1���i�x�ix���\7� ��Kꇥlީ�N�����V�N�-<����D�~�;��'�s?(��%�u6U慲��X�z�XV`q�]7�����)���7O
�d����T3� ��J�(N�ȃR;hM����%p���i4��:����׊Ƒ_�(u�.`�!tB�h�bи9��N;c�1�j�VVI\�L�@g�������I�5L+g>���A�>vj�v�E��ז� ��=~���!�?xKV�bU����W���b�N��Z=�Sb�x�`�j��O�Q���y�<�T�MX�*�]�!&>�^�)�@f������lF�o4[�##�L�N��޲,LD�⠭	Hs\�����\���
@�u:,W��?����t�QJ݊Ĝa���g����m߉9�� Nٍoxj� *�[,���Y�E��Pk�b���Z�Ltq���U�]Q0׈�<A�.�uRcK-OEH�b��S�Aa���Q?�h8�*��%�AV���l�:��O��^W�7q	�EV��@'�Q��K�q\Ͱ��x�G��q-
��(��ܯt>�WE+��|���0+ �w�,(5�^"u`6Lz�,4�J>��ƶ'�
'*�L�!�q���pvI}�t5�6�%�� �>��_�'�eۙ�	Q4�%cOԕ]G�+A�����:jH���x\�2�w+��s��}/ey���)�+�I�&l���Q5����)�b)���}���8�l4��n>�C��	R��])A������_��n�(�����_G��ު�nq�[�(�;���R^��'�8�NX��O3_M[ꋆ��yL����U�Bt޺1x��@!��zy�$Y���jpM�s;N;d�1�n����f��@�����/G8��\G@�c�T*��SB��e���}a0��j�;��3��ڐ�i`
�`GV��_�<Z���i��s/{����1&����=M��īP���Q�Π�|�׻��bϒ(HE����!���{= Ajg6�j͚� &h�{��2ƻ�����6=�-�������1E���2܏X%_z��9A���f��ر3Q�4cA��XR���7����+���H5p������	"�X����r�B�4�pZ�i�i5��0�v~ɮ
|�=|8t�o\y{�2S�$!i�B��f�e6.��u�����G��jF
�{�u�'��~�4%�X���J���`k���|é�β��%Y �%��䀩Qq󱂉��]�ʯ/%�[�.�<S�������^���^]��������l��ט��#�����p�8]ɜ�^e�?<���U���G�:d|�T�������� ��@ܫ�?�,���Uy� ��
�%T��m�-ds`�xX����*��y��:[�Y�R�C�82 ���מ��E�N�����������5��s `��db���OE���C0��l̹%�<.jQŪ�ߨ�]�I�UW�a,����{l���5!��x'�z��(��\��goYf*�j�(
j������km�͇�[0�5�~)HZtǧM�o�f=�ʀ֫�e�eN�,x���"�Vl#Wogf�������{��Z�2�'�S�8P4�4��[uL�*[��Vw���õ���<%KHAJݠ:���!�t�.���c��u�B�ԓ�Ap힙s�'��Cw���Ҥ#%���R�Zt�M�Tv��70"�:�~Ԫny��r�(����Dɘa�|򀷒���hs6��$�g��2X:
�5��{�HJ(5��:�hG���؄��Py���5�L+��&�hG+�h�#���Ad����I?��0ˑ˖A���d�����u��|Kj����H�T|ghIT�w��b {V�eo)��l�&�&Q:�����q��
��G�H�KX>4W��?�Y�r���<��� ˩2������,�c!��e~GO}5�_=�A�$�z[`��$N��w��8��
z4���{�U�C] r�q+�EH!޾��������;A���`���P�B]��|�fր��^��> 	�������p� ��/��]wW�X��P� �r����~O\���Y*`6�U�е�/���n�Y�Rqq��z6�?Q��	��7>ĝT��B��DRW�q27���а�.G�f|0u�i���S�@��e ����F���k�(�Y����U��4�߲>YR^�A����dBM	��v�L�I��F,,F\Wޯ*�f�M���
Ի��2��$%�KI��o��-%�U�[\��k$�K��=G�t� Z�B��˖����5{B��@��'��ɷ`2N+*vk:�/o�~C 	ג/?lWV��V�rjn!ud8!��6�[c& �p'�4^wV��Q�G�2v9J��~d})� Z��>�RBģ�#V��h��$�!1p@g�Tq��g��mj]��FwL\$�e��P���V���%��rl"�L�>NN�%�A�|� ��w7�)K�a�)�����
J9||5k�^M5�z����<](׵����c
�mY��%�o�;����y�jxa^k(m�o�sσ�SH�w���'b!f��7m!՟�*����q1�/*���cn�c5߅{F��W'c��n䰅�wN�ɟX���l�MN�M0r.4��"R��<��k�@���}ZRL>���D�����>�:,1�ѫ~���[���76�M`}�A8���)���V1���x��;Q��c:`��>����Z���&��!����g��*m�u�F^�M�-P��
��)2�:�q�#��'Zv����`�0(�#$eOu*��d�^�Mi�o�Q"�~��5��D����$�(r��Po��Z�Ĳ����˞�Mpm���O#
�qŒgm��y~�.���ba��$/Ӟ����vK�{�QJ�ƙ ��EEb7����2n]a����I8���յ4�{{�P?(j ���a�S�<Љ�����O����t3�MIPq��ʤ���?��+�&J5�^Q��k5��N6�		1ğ��^(P�pt`�lB��&H�DL:�[�IG%0�	A1}�����c�9� Xi�U�%��T�
ucΏ��AY�ů�B&�0q��\�W,��(ts;�>ͫ�lo#�U���`�y��:��M�3eM6{$�]����b���PI�j�=��o���j�XШ�Ã�����C�+�������I-y�`v���=�Z�`�jԲ�"�8��_�\�L��4����)mρY	eR����������q������qq4��:Ʒ�vÁU�i�n�<�G!��sP��hJ�Wb��N\gZ�$0N��&Ġ�Y�ɓ�7V�Y[�7�yNEt砠��Rq�ě��pj����,�]�`������3��b�Zm�+�X�%#~�us��*�N4V���߂�4�5tY��>�q��e��u���fR��x��,�ҧ�Z����ԗ��*�X�ޫ�Q����G��TP�Ad�Y���=��{�'�&�]_wܜ��\�X6)���H����wڻ# ���z�+s�.$���L�f��5V$��ьP7����yo%I���� ��V�!C��Zl)��DG�\�t_�|�_������5��g����}Gx�R���G�D$�*��s���V���:�09�����{S��l��>��Ҥ鬻Lc}-���\�[��<�uM]wZ��Hj���@��:)��G�ij@�Ӻt�4/k���w���0�mϿ�%�L�m��e���kL�%K��M�Cƈ�=�n<՗�(��p�u~�-��q��/Ѡ��W��X����	��,<��.�Պ�����b�+�nA>r�Ǌս��o���M2�����B�GO�Cb�ƥW���\�iA�y�?Az��%�?�c4�����9�C|F�z�)t����`�7ބ*������A��1���%�j��'�V9�����n�"�*�������	)�H�4r� ��r�'�)�;Ѧ��������ͳ(�Ѱ�ܥ��E��ݗX)霁���K��Mr��1�O�3�*p���)<_��Wo{9'�u)���$���Ud'3�Ƈ�*���̯w;���ӝ�,m�������2�p��Wi�j���w~s�� �
t�0]yvIP=���F2_3Ё�5��Й􍾰i����≏F��/�x2O������������d��0P��$��`z%�|Ϝ�˲���&�j��.UX��7'Wq�G��`�����	JSb���4��	KA���?*x!��WH??a�&_� ��8G�m�����:עp~�!�$�t��K��H�|���&�Fi�9-��<Ϸ����<��� nƲY�5����q�:����Z"���K	
�4�_��=�P�S`��s�#f�܆��7�G��!D	l:�c�l_G�T�?ʾ�8��z�����(@���y<����c	4��{��h����}m~W{���S�t�Ad=TB�3}��!B���>
x�*�"�F�a��gc��{>MO!�utdȱ�l����e��y�O��7�!_��KI��9_��Z���~��S[�c>��)��$�� 9,ܦ��$�*���j�D��H�RQ̣91��KKxg�G)��7����wj=Ѹ}�?F�
�`�qI�jl�����`E��]�-�><�;�qܴ
5�Q��ī�=՟�[F`偩>��VY�� ��e�
5�ɤ�-�28db%�vr�@��j��+�$G�7���˖���  w��$S}��d����T�n��C�%��]�!8�L�9�C�(7`����@�N��_�5�J ѡ��]�W(!j 3�d�$hy
E�րe�~d'?0~7�pҒ�NA��B>�`�$z�	�M!����n�+��=�m�����[H��	�*����{�
�~?��)mV��9ߔY�S�#� #j5��Y����"jī���T��a���|^�A�'��^���p�nȈ�TLIX�(_���Rs
[��	(x�M��Ǌ���p"��/�E8_���ɓ�_}áL%i�A`��A��Z�4y�^B҄*�T['F�o�~e8c܅���&�ӝV�K�d��X��BuV�]�'���t��4Š'Ќ�	���d��Ee#���ⱁj41[��.�'��������Yˡ]wU�J�@����q�T��r\�e�0-<w�Ŀ�-�����-ss�7�{����m�幕���s:aak�����{wðs��'�Г~�R�0�g$�9���%�8G­2���{i��ZV�+����h�kT��B���6�����\<u�h�\��O�9��o
LH	������'��a幐irw���(f�XS~����`�m���"�4l��n���)���h(��f��8Ҽ�^�5eq�����uM������2�TT����$r0����\C"�1LS��1����f���E����HӋ����wA��p��3)�<�ڢJvQ`����%1�V��XT�>.�#i�w�֑')p�� �,t�T��+�e�����j4�#G:��D�����y�dQռvD2�y\i)]ޔ���׽�%
/$Zn k�ƣ��fߙT�%��vkI�u�?>��z��yv�l�+�hS�0�n�e��M�h�+�I�n}C�Ŧ�?J�k�< ��4iy��&�����Ч�&�q7�����lx�ǅ�� ��y��H��2�bn�ߤ��+� 8��!ۘhE�B�]r�eh�Nj
�Ʊ�dW�Z���I	����^�L�/�ePpe��58��*r��CÛP&��ݣXv%�m���b����P�r�1��K���\�=�w�k�X$��k�R��Ꮶi��\���n'��	9ʷ���V-vVnVb���f���齒�8Z��L;��T�Aq�L����}Yճǀ ^�\(�^(����YVR���Vux�T�=`�`s=�� /�C�́�:�s�h�B'��L�t۹�P���W_�HII���z L�վ,}���X��)�ߗX˲�J�UB�H�]�!�ӣc-����F+`�k�!D	r��t�*׷���WK-��+�@K�uOS},����6	�R�6�yjL|r!xp�r�wgmc���̩�VW��䅬��k�x���[�7'�߬�dǉԐʒ�+v�}"3b�C�]�K �I�i&�V��>Ӿu�D��N(0��gE��rX��;\yD
h�ꔊ�ة�q�o�l^٘ʢξ+)���L�cn����֕F�zQ���S�U����w��]�p��W��` m�J�3µJ��L�G�*nM�K4�ْt���D[��I�0w�禣}I#�DAb��>E����������8�e�鉹C�5\ŭgY�/���%oK.���od����;�a�}SV]T�N��t���<���!����Ɗ�љ$o��ӌ���ʞ0 c��m��:*�B��/�S_�0s�<�I�hQ����|"�Α��#���.G���\>���U����7���%�Wu��dxs,�DZ��߁�f^6BE�[{CJ֋/�u)Ho�E�R.�y� _��+A�Q��W���"����O-@l�g�{�ߝMI{�����pi�l��X�흂B�48��n���%. 1�z�O�T�o��O�8J��̕Eqy��� J����35�J%�Hgn��\W�uF.R��0��Ѱ]�,N��c�r�-�=���0����0�>�Z���f�ɬD��2�4����1�����8(��K���7+�$)ڕh�G�2�-��%�4l�Rnx,���a{2�0�YS��e�5�S'��D�W�Jw���L�.c��,hPd�n��z����Bf��,>�+5�X�#�q챻~*(��i��z!��w�ifIrT���Sb�STq��I&I�J��K�'��h�&��˘ݞ�0~tW���ZwD���䠽�d�gVU�=�\���A�X���v��_���tx�L mh+���zǲњ��9�PP��f�B�දf�>��ɣ/��A� YE[�i	o��>�+�m�������(�2;����x���'��"z�� Nޛt�q�",�^��-k�n/�i&�֭����~��A�����I'�+�:Gc̴��6��q��N��@�;�G��l�y�U�Ա���n���n|��]F�~������]';��ѩYR�YVg�S-���C�'�9��e��lN���(o^&��o��鬥��3{6Vr�}1co�Tڱ�th�U����f�5�`(UAƍ��%paڵ��1�m�w	���Ȩ�������d�� u��7J+7�b{[9j*@��h������e���#���OE�xy�l���%��<��h�z_����7V�n[*?]�W��)�9kM.�<��@��,�k�1���Ӟ����	��j���0S�9�EF�e�$�H =d����m���v�qG���>�G@5Q}��� �u�dOZa��2���p�����`\8�T�S2���M��F�s�2�8��t����GtrVsW�R����q��M�OW��Ԓ��j雵�����[�vS#��<� }*'A%%ͤ���y�&�k��k�j��W:��Y���y]�cPH�#ѕ~��p�2��j!hަ�A	5kT�'�#�m&y�g+�٧l'}�J����rо��EÅ�H�A�d�au��`�6H��g܆P�Z���-sz�;{� ���d����{�� ���u៯
q0��d(���~������\gMf�V�K�M��0( �Uq4 ?�����b8�k�������n��~�yw�y}�
�N���?D�υrJ�xuj�p|83V�l�J~��/~�ɿ%.���I��g��u��-%��L!�J3<�1w��	�]R��"]�S-��N��rUq��υ�FJ0`#z���N���`��D��B�:�����R��]�ha�8�m��c�iwc#��/N�~��c��%Ѻ���������kB_�\]�QA*_.��|�m3xf�L��e\UO�S^�B�o Z���zP�t�pl7���A��J{ջ΂H*�3�*�'�Gx��ص��d�NCJ�_D��{+��I�@��b��Pco��GPi��紭q�N�a�:F���5xE'n����$4'�CsCB&����?_��c��y:�Q���5�,����i�P��u�x��Vyƛ�O|S?�A�� ��w��(!����*�t�b�^��ـRM�K�˽!11�ޯ�9N���2FA�Puۙױ%_����P�s#�xk�2ze���aDݻ�;�P
�-L{a�YV1U��ڱː��܌-�&^��϶�C�-h!v�z�/۫��:�e�������m[�嚿�ן6^2���� -9��)avI���G/�߬�M,%��x0�7�1�l�����lе�:J�A���Nb._��U��8/�˺�,bȭ�q	V�4eM�v��By�C`�ڨȓ�BK��'��+��X?Ph""�����0#,�x��4=���¾6�V�
z���M��}��P&��H�:���G��\��\��a���\�~�0��%��U�4���wX7͎�	��@���P��gYx�m�p�m�}���ДI<�K��g��^1��=�����a����?���ͼ�ł�y5�+���GT�!`�SufO�h+���O�,\q 0�ߧ�(�4-"����U,�c�����QsɡbU�1�,���+1��"$�0�l���
q�*����9@����U�ߓ�S>ڒ��ٷ#�D�sD�jO��cF�)Ie
o��$V��9�klt��-�1�fʈ��CUj����#F�Y��u�;-��O�+y��z_�;I���I����F`�c�ѹފ���=�|Aa�K�b�x�ɢ@�Ĵ�����0�s0Ά?O��YA2m�V������N.�Օ	�6}����h�h	�U��,q�1�w�i{�<5[���9u�TR���U��q�'H�ȿt,����%����H�o<Q1�o���u����x�7������J�W��Y����P�!I�hrҜFH7_�>݋qK$W����a��`��kV����s3}y|c��ti=��ˢ�UR����bĵ�8����, ?�[�Q�Ge,�*2��ޣ��m���Q\��7�qi|d��������vWOS%��h�_���>.h�,��N�)?��D-���O�
��t��S+�N�5?]��L0�.,I��4��"U�e7���VaY�if���CL��q��;aЦ[Q� �M��{2���6�]��iA�	wm��`8NtZ!6�}�D$c�D����Z�˞�f��t�]|��%�����8��}�7^�$t܉�4Z����Ze�m��BH����$s���g���	K�=��	c�y\}�_Ɵ���aaR6_14{� �	#>�K�������a�<�G���_E��0������ބP��8-4 #�*P�ԧ�]@?w�Q�q�g��4�D��f��3��/�)+,�g]?�D<�?����4�i�
�z��6�9�Zd}��SA���TT����/�p�̒�ܔK�p8���<�4����3��Iv�jt���k�/0�����}��}7ױO�������m�ߘ�R���c�Y!TCP���^������]�Y�^��b�/�
�s�g����=���T��5uw뫋��L?] �*x�c+P0!*���栯�Q�r"�����d��%僂��i�$# ���"�FjF<<�ءZ������� |�LB����"�yNv�1��:�N�h�X�u�G4k�����׊�\4?��O���=�($��Ʀ �@:<�\��1" ���n�^�q'0j��o=s֧Z�`�a�q��'k��Վ5��'S��m��k��b»VU%;�lv����T$��#"��C>�T�q'/o��7�y9��){����S��Q�zG�b��{�h� F�l2v�`(���Ӗ���
�3����\T%����Oo�
�T��{�(��-D���EP~C%<}��{�\��`{<�ULu]���:��@�)�?��۟�;��@@�IE�����舆�˱��5�3^მ����+��'����Ю���g)4��&Q�AI~SD��_#����*8$l���}�(�K���\��Ė�����qWՆ��Z��7c2���f���|Z��t�m&�h��p�9�- �^�"G��,$�H���b�@���H��^���IE�cmI��s��cW˂����D�ۦ~�?'�I�'H�����;y��g�Ny�+�֤oTy
��*���U�B �1|ިl��Z�Sa�[�[�%�|{��W��`� M���s�S#�^��;Ι�O��<�h �c��}�"��O�+s5A�e��-=�i��d�l�׭�c���>�i����ɯ���m�ؐ۲��gR@Mݫ{���������ha�6*�)ƞ��u~C�?���z�=��^^�|������椱��HC|���s��i��QX.T�6W�~�"�	<�8�/\
�H,� ��7�X�llj��$[qY���9�%�J2K�dU�F�z�<D�թ��t����(��$�z�j�B=�_�q�O։?d��C�ؽ�޷(�a�)ɧTS5||ܟr�0�nO�Ymy�NU��U(�\�NՋ�Tow�9��Fz�]����"Y�T>�)f����ٸ�E���}�S���nL��t�t~�⭠��p���z�;b�J�)�Ր����䆢�K0� y%� ַ��&���������Y�7�!6 [Kݙ��p���W�,�|H��@#ӳ/�S�4֝�����t !�oYt��5���EG=�w�4���=3���X�QɆ�rI�q+���ҶCb�?ZR
�Iʹ��(��D;?�y��rg��.�Z^�a&s))��[ê�T��R����<��{Xn��%@�F����r�����C)����֪)j~8I^�MЄ�ݝ�)�
�;z칔�eR���o�� ���qf;�ٓ�
�m$k�	O�����{]�7�i=��q���+�Uv����@[