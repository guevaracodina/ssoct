��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ��p"���C��T�fX��k�+��)��6�'�3��$���)��2�+�
�#�7��Ib����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��p�@n��7E����������kи>de����h;�3�������=���x"N�X���|@K�������1� �!D�L�{N'�u�C�4OeՄ��vy�>Dl�H�T�����T�h� �~OM*E��CJ��#ڇ�Ʈ�pB�����"U��/�7��T�K�f�_�0l�8�����+׭�͉���k���F��i,L<\S�� p� ��I� �ӿûd�Ϛ�kB�~wB�t�'�X�7�w��EO��?���*�)�W������z���ɉ�2ft�Uk��5�&�>!��5R�C�n���>^��j=^����u)�Æ��-~fv|*�����T.�n�m|8Q��Yt��A�s�]�g5)�"�!1;Ʊ륰��P3���XT6����2�
�_CT!g��.f�
�[Y@h|WgY�P��y\�� ���إ��X�6���ܫk֬%~)Yhd�	R#=P�qp|�D��t+���n&Y�r���n��E�MA�t�n7>�W�Di�Z'�x=�(��"���j!�FkptA;c���D?,cz$"c|_�5��dm3��N�����o'�π^��s�[�����E�n��m�|*]�-pK ���1����9�'1�P�.:-��WU�e��"�uI
h�h�O�����&|M�ZML"��y9�3�F��s�3�'#?u�j��B����ţc.t,v���Z��c`�F<.��R�j�}<�ө���mA�Z!z M�o��$����l���8�yk������_�ɇ�A��+�ܜ���M>2�	�
�5S,w��K�J&a�1�l�j������^�ܧ%�&]��Qbx��Fw�)���C��#��W��p�������0��:���q� uK-}���}3p7$p�� h�"
����M�E��-�A���N���%��J��p�8O[-]dD��Ǟ�b&�� b]4j���̬�*���Pj������U�	H�L+{n��;O�=���.G�����jZ�[V�e�Aπ��Q3ٮˇ>���R���rZ�-"2/�j1�Gi窪�g���iC^�"d��7p�n�d��h��CA��������>ڳ/��F�U/4�n����1�~m4eɴ�{�!�Ăd�)��g'�y���6�i�@e����U�����e���kY����V�($ ��73���9�=�:���{z��o�)���X���L*W�f]�WA�1���������-����R�i?1 (�Fp���7ؠ�y��
]׺)��6������{̋�N����
�<|����2&�����8iO����`���6^�JKqf-��K9-4�+R�c�4Ŵ��zo��A���n˜l���~AYۚ}06g�Ȟh���<uW��XK�.���S���rB(��ٹ�6A+pќ�+�
� -v���N��ԝ5��]~O��$��a�t^uB-ܧ�l����?9�ceS�}��4�0�7����1;[�`_7�#ә@0P|�D�����*����/��-ν!���	�?b`�ͻ�u`Q�1V3�8�_��	��,д=��]�h�[J7�!�;���>��s�m.��|�#H}�1�Ú͆��-�;�����_�����d �@i�O�?��x9���(%DJ>��R�����s����\=�^�f̂���U4�yչ.Yh�"���~c�L,���z^��bMg�q�t�^ׇ���U�|B��߼��.�v�8��B٘�#�2!7�_%j3�2��h�TcN��)*��,�HR,`�l�B|�2��_,�f�&F��|��WT�=u��I�|�S���i�VV�`�0�M\�cT$�S�����v�f��j�d`G����$o��y����8Cj�,=G���?��ƸX�NJ�R��:QR����ǉ��#z#v��W�Mĳij�v�_�B��*�b+Y�ݞ�r�CN\M�b�"D.��A%-;<Wr�i�M�Q-9䬃�Q�+ń����l��bE�C*�|Ja����
�C���Q��yw��ԡYxD8�8:C�:�!mI�LS���4C�R��2}�QI�ep ø/>�T�$��ǋIS��Ӻ0����,�������<��B�\�I4t5N7���q�\����lD9�/�b-�b2�eR(�(3|S�Ĩ��W�o�pG�V�����r�!&�k���K7�l�g���>o]ˮ��ޱSZ-ĩǷ�Mp����\���B������^>Q0j:�?�z�Qp�o>(�a,� -3�#r���񞛝;3�n��ϹS�DV�N��R���+��,�I{������].�U���;@o��>��$Z6p�[ȭ�{�g{�uN4Aov�W� \1��W�����w�Pp����nA	���X��d\+�O�}�vFر�����D||=8�f%��0�%q;ġ�C����#|Y^�	3L�������[�L����8z�Dg(��M�޻2BAG�����?iB8-�������������g=W��X�g=zB�Bi�+�)$$g�L<"(�1��R��T 8�ޟW��Ù�%���C���{�[֫�BiZ��}�_M)��0�{`�l��\I��&�Fl����s�ò+2	�lۧ8D���&��������`�y�Ȕ��;���6Z��m����>x� Wȼ�U��ٿ��4ህ�}s5�r��U�ݽ�ATB�"�p���^�`�&�QcT��M9�C� ��0�_j,?�'F^�g�6�Zt��љ>������%��?2Y]iaBy����*�"��HC<���f9�I_�*\� gAz]f��B�'�j��?u�r�	�jY�9,~ܾ��_�A��4��I��ZZ�ld�Zrn�W�,�*�@��ߋ�_<��=b̯���0�m79���]���6�Ǿ��"&�4ڡ~p�Ւ.B�A���7��d��)z ��`7}��9���H����T ��0�0y0��^�I0N����>��F=��7�p�)<)g��<�B��ʌț�R���H�m!b��n1O��z�V�a��xL��.8q	&�iVX;}K����iv���0ٞ�U�d0;VT���-hH!����s�j]�ak���Q�#��a��$�~�A�H��g�pFITx�Er���kЇ�Y�Ȓ� �Q$J���aU\n)c^*|�;