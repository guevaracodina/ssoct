��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ��p"���C��T�fX��k�+��)��6�'�3��$���)��2�+�
�#�7��Ib����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\n��a���5,�dC���
��E��ɳv���3�SX�v�P�-ѺR�1��БdZ>���>��AZ��P.G}�3�.�O/a�
��Ө��P'�Cu;tk�4�χpt����w��zҤ���4Z���="�U����ᑠP�S`��1s�,fV�弨N�՗n �
�j�Y�1n�ǖy��3�Hu}�_��O��.\S}����f��A]�9��w"�ȸ��4��/O�7��Y������n�k\�O����� X W���#��t�-f�s���>�$�n�͘K�l��:�|{1W�2fT}(az0�1�z7Ո�bi�
��U����#�!�����2�j#��TM��r`VP���њν�����<%K{N[��	��l������N� 5RR�PJm�Sf>���x6�-��qǍ�B�q�9����z��ڋG&>�F+�ߋʛ;�LC1�{bc��h�n�~���P%���'@�X9�Σ��7a1Q=�CC1]Λ�J����l�W�Z�c�z��1,�D���[�zN�n��&ɑ�J�]��5F��1���W:!%a���JJ�B&�J sTA��w�g��{]Ɩ�G*��h�y��4���^M�/�1�}��W���b��(!㥻�M8u}�Jϯk�O��i4RBƤG�?ƺ�����d�R�iWC�Xx��H-��2mտ6���"7�^�:����ʐH����\3.�Lb��1���R�Oc�HD��ƨ��D�<� ǝ1���B����(��ãF��1�M�\F��r�BT��4Qנ�7Xa9�D�&�M9�@=������ɂ�f~V��@�Y]�o�ʫW��]��v��
���6������L]Y3���������&B�o��U҂�P+u�|m��W������1d�t���F�8zՁEi��{e�,Ȋ��k��!����}�;�^��:F��5�D Pj���;\�H@: 3��)\u���P�#����t�p	=��HE� �h���h�v��o�d�f����^9�M5�o��3��������4`�w&�(���VY��>�+]z~��X¿3H��T�n�n5jF}�j���#�^w#��p/KL`Җ��7�&��/OM��C�
p�/���d���~��VRU���U�ϗ��3��	�9��uL��.���Y�"Av#,}�������dL��U��Ϣ,	6+.��N�re�]r���U$b4䯡�M����%WdS��\�2��#'��kO���Cc�a�9^�h�?va��-����e-D Ҹ`�0�B�O��\ZW0a8NP�q]L����d{�H
�Z̯�_:W�Z0@��o7��6"��E���v|?�]TD��Cg���ӻV�rl��5O���W�zE���M켙�LAZf�%$�)�j�f��d�|.e�`��x��r܏�K$E��܏ȭWoY�s8�2��3����:��_G"*V�/к�И��H|@�	vu�����s��0i�-�������sx�JsO�.4�D���fw�m�&�̤��y{�Z�G$�2���
F �g�߳؍4n�J3
�����g�z�sM��y{|*���#�j������8���zvꒈ�9$��*RX�_Rλ�y��F���l�D9�~`Cn��K �0�7^���@�ЂBǂR�|UC���gt3�6��wZ����	�/�l�P�Q>s@�bah�$;c���h�[Kt�M̄����O��5lD�u�D|��$)�,g�!��֬-��E6_�,u�'��2�k�1� �_[����iU4!v�L1 \{]sj���+h�ګ��n���B�����~�~�%�����[Gۍ�-�6��{��l$Si��:��U׏������U�5�5o�������"S��\]e�b�vgb��1:T�����	�"z�C�x�_�c��S�����p@�#���n�������9D��ٲ���q sp��܄<s��;x(:�\��Ďę�U����Í*��J\��ڞ�����y���1��S�z��sD��K�؎'Lm3Ȧ��mR,�tي	���O��u��`�+�v]�wǘ��1�#h��]��B��\��}M�T@m�"�[MK�8��țA$β����S��m��o���#i.z��;�=�p�� �
���>u�H0D����h�w��S����,���sW%UŃ>�x�B}T�'|�d����T�k�ڡ�0������a��<���2[jH�]�������l��wL3��O�@�X�R%��a?�	�+����gai���W��=ۯ���nA��uݜ��❩�z�ih�̙���7���q�#�"4�]ʵl嵫�����ZdMH�v�b+�5�M��G��a�]�%�DG�j�;K���K[�绯��EV�+%�G���Ԛ�^��ѐF�I���6���7u0�C#�[������z�E��k�c�:5����A��&dW��E��JkkyDo���*��(��;<�KO���8�����>-E��Os�:��JhL�>")��~x���or��TE�u����`	l@�9�o-�iUYN�sr��&�w1��S�]�D�Ε�t���y�Ĥ�Μ���Q�Ŗc�ģ�4G#CI)��A�}����c�k��4��t�D���P!ö�S<-�� �&Qk�^�5tr�:������w`m'9å��1���sKx�M�Z�.��	F���8����5�����V){B�$�}�bLv6���������@��Q���0|2�W$�Z�����T������Wǘ��Ͻ0x�G��;��Q�����&�ޖ�1k`�I��<s���Y��e�����B�r�F���� �M�S9HL�M+�4w��������ݼ :(J�P�9oV� ��k'����_&�OjǍ'>���s5�ԯ9),q��C\���ʣ��Z&��VK�a47:���[����l��7�ls�4I B�W�{.��H��v1W�}�C� Į�@A�Q�PDO�#�&,��
�:���􉼿�><�z���=��ge޳`(6�,{�VDJ�4O���;��1�O�`Nq�ї/��284�c,b������A�}��U��|�8��ְ��4�����&���ĖXP	ß���P����6��'�����(�������u��V����z�0�C�ⶇ�k���]30���$D�����_S�����G�&����[�%  ����s�w��}�s�y��@]dx���0!�&�����c�3}`椯��! N�O��*���$��v��o�\	al���u���݈��P�x�YQ��Q�)�U�7��K;�7��1�����{�V?��W�NȢ�B/h�/}M�K#H`E�%㣰�p���W�!�tB�m��܃g	�5��U��>j�S��>Ǐ��VU�Eu�u���w&f�;�Ù�r>�\)�W��~����l[�-�­D�T-��^<�K�1�w�_��<�~⪣��upC~�yg�8���'T�/F	�4�HidhI���4�*�����P�3�:�Ԁ�]A�$[�l� �Z�?a���pAx�=ݨQ��`�Җ��Gy���e�X����O��^�mH���Q<�Q�������9��g�/���/��o�9�*���p��=�/y n�{{g\�?�$m���e`�Æ�\()ZE�i���9��uS�ɘ���E����W���7J�]�T}I�	��O�9�H��H�����*��*t ������|��G�p�,����7ƾ������j�W���0��^34{e�r<��>�%^S��/��,���&p)��)b\e�2�r�8�1+������p��C1l.�@Jvo9y�Q��R���R���G1@Q`�3[PA!��t����֕��	i��+��>�ȑcᣵ�/�2ԧ���v�R3���y�s��r�-����W��|Av�-��
⺎iƼ��g�i������2[�tFz!��
h˛
|ʜ��mY�������R_�̾�	����0��wZ�tӱ�*�!�Eknu��s����R���b'�}����d�����bSE��s<y���ld���.���y_]D�>�uʧr����4M��A�O]ȷ���R��m���.Q~����Y7?7n�h�WV���K�.ӎ�\>�U\�Z|ī	���.ƚ��� Q����([0��4q��\��!�����&O��`Z=����D'�t&bf��"2�O�,����5��d�:SKg��VZ#v��ౄj��N4��!�Hd��`�x��L̉q[��bR����
�����;�B����ísԡr�^u��fad'�F�n�%k�&1�7�n���)H���j�N"ob�ݚӲ;��&w��t��a����!�{:��1o@�Q��D�XI'o���O1�x̊2[n��]n�B����6���pĺ��!kKd�DsI�����x�#W&���M�U�ڷ�鉨��~4S�Ե�5�FM�m9+�e�;߬�}dX���\�&<P����]�\��ec��yf��쩑�9�ki5Ƃ��K`bl�\H� ̷PT��`�pX��|ؖ"=Bе��Uax��mSW}/v�c��Fz(J/� �����v�(K����j��p���t�zW�7fV����½1̄`���P4��_�?�Lxi���︝���)��-wZM��3�T���V�4b[&���!�Y�nb|�#���֓��fo2( 5�E�/N����ߗW��vs>>.
`�;��g�oix�\�7�N��O|�d$7�k�\����ڣ�����j����I�Tiaf(�~�(uʣ/<f� ���2u|�+�ݯ1�ֺ�K�����ϒ0�;xBS�O:ϓƗ���ݓ�oY�c�}\�����;�m��#\,+��ϯՠ��I���Z�O��1�����pt�JK���>��=�v��l�S\:� [~"v�h^ʮ'���9ld��\�I��ξnG��~#�jTl��������ڼ�W��7||@��Λ��o��PU Ge��K}R
�B,��T�p��ʍO+
�f3�_��Tl�O�9{3�}�O�7t��X�x�~H�`�	v!�W�ɐ�o���X�r�#ƥ��a�Y�8|��-f����X�"��?	!J�.������k���x��>�Ԏ`��s�l"���Ey*��J5N�'�n��]�T�{�3�da 3j6��S�`��ZK �6�����	V��Et�G}�Y �j�D��N1��Zi6��t�����,�}�{ڽ�wX=�˾�߄��ql���looh!|1d3��D1�;��@����j��T��B	�L���y���\S}�W*��xq���g�,7����C�V�1�|v'��.^�'m#E�6_�g	 i��ua��v�MIa����O&������m�F3-�K�x��u)k��U���9L��1�
�(!�f�/� l}$sL¼�Z���Y߮f}|u���(�H�Azm	���se�,!}JiG��$p�|�~��<�;��Ko�K�9{ے��������$W2(����#��^��،�����>�Dm��r����]�n�|�_���%�y�B�0��E���������:�g� �h��^��?P�iD}�6%�=��z �- �z���Eg��j�7q����kz�O�ɭ��Uط����q4k�l�`hQ�ؔĪ(;�E�1�kr\������* ��|��n�@	3k�̦o��iH���_I�b��C���Q�cK �����k>s����0L`I�-���O�����d4�d5 "@��S�;T�f�MX������ѳ��!;p�<��eW��C��Ki5�أ��5C�o�8{�}��{vY�_E���]����M0�8>��^~�4�	�0 f��<�䒶ͨ����\ă-V�|+����~ �Az��N&9^ߤH�(��#���12~�i��d�6�4\�VA����T�j�Z���5�i�#I�RU���_D���e��jK�-W�ЍR���}��}"4�i�y�ۈt7���nu�˺K`%!�E�I&n��9b�1p�!r�8=��sq/��l��._�!�z��p�	a���̰a_~�2���ExN�Z�}޺�'����,�Me3#��k�pKp!�)_�8�[d�wi�,��*���}��	�	{�(��n`K�K�31���"��$.��?U �X�n߈2�pf��}����Mu
<Ie���IR�T���	_�'mQ��p�hi*w��+�c%�{sl��D�ߑ����	X?��m#P:��=�T{��]-��an�g��brT��}L�M>!	�s,��f�ob��h�Y���>�����FM�Vj2\[��i2l1T�
di'��♧�a{��,�밙�u�pʚ�v�c1��(��}h�?�n�(�I꘺O���Ԁ N����F�B�$d٠�bā�֛��*�:V�1�J�<���_�O����?+�<������@���o��]��OcC��?A�	�AG/���M�3|�R�G�9��?���8�pKDc4w�$��>70lc�ګ�<l27���3��h�mę����ǌ[c�8��Rg���l�s�P:Q|ke�W��@h1�����@ی��N��m�>�aZK���6S.��9s�:C"mi)����5��̟�rҐ�o���r��z�6�����������A��@����\�cKY�F=Yt�5O����Y7I��֝A�(88�Wך�v�^��JH(ń����ɳ;�K6u���"M&���&��Mt��&P������#R�w}�3H���M�_U�7����$1ϋ�;i[t)F���=wA��A�q��c�(�`u���[�t��#=�<���^�6`�l�V�
sԄcX��2׏��=�GAO��@�Sة���uC�XF��Q	�ٰh�:$4�@!� �/E��.���j��C�~� v�q��<!T��f�Ԏ6��6�?���śθ(��i_VA�"Ʉ�F�mj���[�a�aTu��SKdoS;��/a���b�U�VYk�ߏy�z��+1���
�����gA��\\�W���@`�ag��("f������@�N�(���#���.�H��u��x-���[#}�{�z~�I��j:s7�~�m��Gf���^|9��Ƨ��>"��vD"'���a�a!�����h���t���ˤk=+Nl��L@\�'�)�gk#�v�9�w�?j-���񵽏w���Gmb��f��X�lI�$[4�8�η��V^�ּ\�6��A����r���Ɋ�]�ٮCj�(0�l�&�\�P�t��eH���q6
�b���Y��+�4x���#м&���s���\H[�D��RT���y�joӽ�yQ�v�}�e��g�DJ���\��+'2ٸ��7 �����1+��'����L��]�Yژ�W`����v����N|aV|m҇i�����T�Z��E9�ڨ��o��cs#��u�}�1k��L�y��I�x�������5��TĄ��WӀRj��z��%(뿫�w�?�S^@(�c̟4 �\_�ܱ�LŽ����!�T<_�	1SU>q5�	Ow?u� u簰�'��{R�C%|�~���� &�p�Nr�MUNd_���k,�g�q]�����D�m�Y��g|�r���+O�'لf�j�q���+|���rљ��H���={�����d���K�'T�U�ocM�ۏ��
	�) yN}#�{; �wkE#�mI�u6�7]gZ_�~2\� l/�-�&�E������K�h0�%��w�z 7ї]1$n��(-�T���� �;!�g���$V�����P%Z�ܺ5�u�o�$5�` �dMӼ��`K��p��^�R1S'�X�L6#L�b̐�D�髈�>��;��ݟ�9�	eĪ�|�p.���
�A�C~@t�X(���}0�NPr�ܹ�
f��\ԯ�aÕ��<�Rs�7�������5k�/{��J/`^S�-�E�X4�y�������4�5�|��l����w���Q���#�!]�+g�OܕKy���ߍ�%�[�i�pr_@��g7��"��^���n褽U��I�h8�b�v:S���s�������P��vIe�*ߪ#������]�3�C���9�����9;}q!�v-Aq=~(́7�mT�3� ��l/kW��$��������0E��d���Oy{l�o4���D�গ�&%�$����U�Wp	Yc� �:�q`�1 ��sq1���+56fsd�[����|�l������q���и�b���� >�U��MM����!�k�3�Q��� ��3-Tbh���i�{oftӱ߼�u�+�;��ϾS4w�=X���B��c[�1��)<��~Ca��X��L*�Qo`��1"��U 6!P�T��_���Ŕ|�C������)����i��4��ױ���(�b�d�#�k��D�Av���~ή���*�����>Q*~��B)��@�o�"�2�F�i�\�(���v�	�֗��v3�dս�oF��k�EVp���^�6ew�.�=Uwph� ����0M���㟛\��@L1_h�-9h��bjv��(֦��OiAF�-pp��q����1��Y� �}��UX�����R��Q���+�!���2��~���i�|����˻"д��P�'��S�S�2y\5�y:N��������h��lY���K��i�3��~G��{�"WL����}�a��.�|�F�D��`Z����l����@�j�����c�n��`��UDW��Ă��}��o¦n���$E�j>�}2pXc�j�p���m�W����y+F�kO\�}܈@}�_�����f�MPN���FJϥ���^{��_b��{R�T8����b�K��\��Mz�F�n�m'���5��x�=���y�[d4��0��$M�r+ws�Ħ��F�Z������I+��h�x��z�a(T�G���T�@��h�f��e}3FyH�ϴ��P�ǳ�h�< ��#k���z��)^O�S�D�3��5�3�N���o-����%��+8j@(:Ej���̘�u�k�g���MQ4mi���p�B��~v���Ė�+جW���]xd���+�� �O��r�\�ʂ��'U7
��r�g<��P��Vs����	�
C)��UWN�嬵;&��y��(��ј�0�:���,0��\���s������,Wl_툡 ����'Am'��JcbG5W�xླྀQ�	��cS6�אhzk��=�ʗ��D���3 ��~��Br�I�a�D�A����Q��$�:�9�����X��@���qR)Q�LO�9X<�a�b�ǯ�g�||�ڽ P}�H�%�X*e���!�<G��:�J`v��*J�qmcm����[�D-���7İ5M�x�ԧC��qg�N��\9U9-P�(�雡nf՗d���(bV��$�3�!LT�*MFfa���ڌ��{�g�AzoV��<L�����v�TN@�xv2��M!�}E�E��] ���l����3�ի��U:����s�G����s_.'�:u��� �+���Fr$�3���ڛc��� �J��
-lL��&�$80*���uձ�]�E�� Qb�UO�q}���� ;}�KweU}u�<��y�X:��U���������A���;���ʐ�v�/C����)Y��(H��Q�l; 29�`��J�7Tv�Mk��T��%�}s�]g��+j�8�"F��Ï�t(53�s�=�M�2����5�-"�Fz���gH���v���:�!��>6�sp��X[)=yy�~��{#Q�=�Hx{��˿p���=k�Rc�mY��w��%!)�Y�u�󔓡l!a:^��Į0�/�3��x|����hҲ@TSm#�o$���_j� #Xk��2�s���VPQVH
d�&m���q;����g����Dv5(TI��i���7A�ӯSݕ������ei�H����>\��&_��\Fw�3��NF����l���8y���v�$�� φ�*ɽq��6���7�v� m�$d�(AV��
�~��ŏ�w����3}Y�B�O"���J[�W�
��y��[�_/���a�h�&2�-�y��$�|Hy��4����9�x:�`�N�B�b@�d�)\��;3|�̠"�@TN��2�/�Z��B�CP��:G���

k���!B\GKl^�C���6-F���i�Y�
=�F�E��#���i*�/�KtycEI�=�b���0�S��33O���<���4vnN���!��+w�,s�9� �'��6l��GK<
�&�У0aR�)�,��D�Oe���g#��J����{�C�t*b^��D]i^��P��(�d�[~2�{��9d��!���_��Ȧ��}%@X�Jt��@o3p)-;ݰ�	mVo�rɽ���� �u�#"e�O�q*C�3F�T������B�+f��}��Ef�j���������qs F#a��}�W��F~���n�.8Jr�R�sw&Z�ϰ	�Q���H�y � �
�\���ȬG6��r��66��v`1q�r���k+e%��(k�ʟ�ΎE��:��oG@qWk2��c�a���{le��{<c���NA[a���~�X�|m�֋9֯��4"��1�8�Y]cE�"/�|{�z{s�͞��	�͈�a�s��Z�nS`k�j	�ל:�D�@�?�f��t��r~��;�5�`��1�ԓ&���Ij�g��d1��8PT�[M��(��B�W�ਞA>?ZA���'��/���w��I�p��4��Zy/�G��c=�H����Q�Q�'Y�ؘ�� $!/-
������68=���I�S4zJ�;� ~���)>��^ﵮ�37(���`.��M8{p|W�����b�*"��q���6��L#X%�ݐ���NC'��
4'�~���LGɛ{��m��\�bP�۷eM�� �l����^Y�|�O���?^�\u�ͮ��'.��y͂�T�xe�1˖f�Z>φ+���KK]B�<'��EFN+�`���7���u�
��+��]h�2�2ِuI��.�2/f�����KO�_���Lo��{��|x�A�,�A��>�@��m>s�lY�Xes�{%�q��FM��[�� �kp6F�2�žv/eR�������jH]8F>�.�՝k�K�Њ@�un��fo@t�a�	�3i��;���;	���(�I��}�"�p��J�$����O�J6����_&N�Y��nd�y�t�ý�W���Qۈ��HC�T��4!��qg��Z�/\�|(�~l����_&W`�	n��%8B�Ǻ�R�ڲ�ߒwi��h}N�g[�Ъ��8Yu0lݩ�&n���#ű��i��R�j��� �g����v�o/���4�H����?��A�ٴ�nX}�e2.'I�	+e�T�֝�6�%'fv����	l,'ԓ�M��bѸ%[H�t@�FG%��P-+�Ə���JJ!sEި�e�V��PK/Ad�ي��r��)'Clȝˣ�A�������%�2�8�����|�iM� #��R����Ǿ��H�����h�c�D�<n�3�_�������k@����4�"!0'DA[�TϮ��}��9����BekH�^Z��o4���`\�B����`�ul�R�Z�9S�O����
p���[S��)�$���<c2�Rw ��*lD1�!q���Oa��`�]�e/h��;+}S�^y/b�gX�H�ަA�$Qj�3��M89DI�L#����:���H+�������|�2�jOn�e�V'YLs�;]�;n]�KXm���5BQ|(t���G�	�
�d�A���&8/�_��P�7		��x{���ND���e�R���f���@D����|AjN(�.a�v;-�s4�6٦�DE�"V8�XK)ONY��7�#�г�E{���7:���D���<sg��?w\�r����,�)�}�o��mQ\`	�S!���A
��G��}W���s��ES�98��P��k>,#�6�l��r}xϩ~t�6�g�jL
l�.v�?�U�#~���G`�e"���]�J��(>2�i��yA�X�i������ ����q�P<��yo~Ek$���*<q���p�-8x ��Y'%O�u�ԭ+����������p��45�M��C��RR%�W��	>�0_%(�nV��Lqx�_%x��o����a]Ы�'8Su-��7CS���t��dK�䗒th�j**V�FyS\Á_K�C�N�(�u,`�%�;��{P�a�m�H{�n��~�W܂���7放���.;��jT4ĭ���u��~�N� |?�������Bz���a�Ro5e�y��vw�P/]2z��g�����w�e�`1�����^��1/V=1���[���2��=��fX;P`�G�~}\vG��d!Bdx�
E�'FjD�|5#�)��mV&J��D�� >�y�M�����]��cӻG::�Sc@�&�mr�o�� �`�?U�P�e����4�-r ��.�8VЙ����M��Af��7�jb6a���o�s�o�����;�V��2��JC���`��Q-'�'��"���]�)PR���8:/L%I�K�����䏭�j��h�L�k�&_�5/���}RBN{39</���떰�_4�ڼ�eM�m�����ͽ}��Ņ���ɹ0�CZȗ�0��k�J0�6�I��O5 ��X�2���푭��>��NK2m���֡b���?�u��Zg�/6��O��>��D��$�I�y�����,��M��[�ǭ�8Ln�\�b�����6�T��~�]�	� sOz�-[�䈨H=Ē�¦h��!>*�,�J�[�@�����]���5����p-����(�����yK6�]T�'Ǎ���α�
ںՑ|�\�V�!��*���@�F1�<y�H	Q��e���h>`����ϒ�	��S����_��5��?j�o�CzN���Iހ��Z�D�WK+u�8K�`Y⋻���N�y>D�Yt�z�,�(��j��J�5
�	��uǿ4��f$?��B�:���r����mO���6�"p벉/Zdn^��^� 7��N�e����2Ӂ.l'�W�Duj�5�m��(�B��h���q+h���+����\�+͚�Q4Cގ�\����R��t�0p��~�e|6�&���҈��}�;�J?��Z��� �=�0�����x@�ؠG*'�tR��eۙm{���X|��J5y]�H��WC����ٴ�`2�_-~��Ԙ��$A�b��� &�)�dF_},��
p�a�Pyz���w<�Ѝ����l:7b[e�_ń~|�rW�+�dR�xiA^&i�d���ڥ	V�M��-~,ȉz�{z��+:BW^V�9U��6
M����{a����9��Ih�Bam=6B��/���n:�������%O�D���a,z�Ex�2A�ba���;�Ѥq�MԈ��DV�0c�Tb���b�~>���˗�B�s#Z�}�S�V:�v�R��}�'��A�M�}�b=�Z�"OxAXs��� ���� )�"z̏3�c�|y
V���[mj��>���ł<�+�L/�v�3��B���y nC�7��VO��\�=	Y�A��
�/s�0�`{�l�g�q�5H^� ��s�����7��_��&���3zl�7�ŗ���sY�<hˣ(2��%8�<�lȵ�#�%eã�w9�kē�W_vax����f�� �F�ĴsQ����ܣz����A�,Sv�_��#���MVRl���N�K�]����$<;�B�K��v�<%�� �ƜJ���U�3��W����@�"$sfؒ�,��96rp�F�b�m��s�B����A���j9s�58%;�~�e���О��������_u����]��]�%������i�!zc.뀴O�ȃ̜M��i6S`�Kw�=��(}�JF��zP[�B�b�c���o�M�f0���- }�+��u���2٩ű�͑57v����X�j7�i��6D^�Ͱ�!�8K�+�;8�Ks���z���+SmF��(��j���(��8��1�J)�|Ǵ�d��Q%�zzz�}�wd�s��|�`�^�NY]$�pU���du�P*��(9٘F!���<��t�w�-��z�XC�6��R�*���m�[��o�Y��F�G�_���z 3:��^�L��'�T�JHo�裞�J4�u�k,'�a]���v����B��Y?w%�����6Pge�Ȕ=�]�8-_�L�jY��J�JW0o�:�=�V�\	�j���@��$�垨m�<)�v��^��
Ǖ�ˌ��_\�������4�[4Z�Y^p�E��(�����rEd�q)#�P��2`6�EK~W�my>TG)�n���䨷�*��"O@�'\��P[���d|d��^��t���Ĵ*��PAf����%ɇ	_c�m��e���>���[0�,�H�E��\
�Δt��6�-�k
э��)��j���noG	HӋ�F5E �|����`�
 ���C�ź����2�c�(+��7��u�-�&��,��V����?Y �פ���:ˎ�a�.[��� �?��G�$��9x�SMymMDAk�ܷ�l>�d�!��֝lPF�V����v�q�E�)D{~2�PJ?2�@�T��j]n��O*���ܞ�r&T�!�XA�!�Jc�	J�N����Em	��H�U��t���e�وO�O��H_�5���J:��B\;��W����h��	_����+H��]d}�"Zl�|��,_�d�ɍ��v�3q�k�"L>�V~׋�:���������	��`'����:�X��HY�ɹl'�� ǁS)(��{�K6ͥ�t@��	���(<r�#��s�c��
�P{	0 ���/dW�����4�OB�&b8�p�DO���&
7ܩӃ��F�W2��k~�iM����ɵ�Tr��ʪqR��WT%��,����]�ϸd�*��R\�W�6�W���@�N:lz:��'���$'<$b<��s�r\k4[��|Á��F��%$��x6v�h[�!_�ķ�j��q`T+��e@(a��8x�R�ۘ1	��)�^��@��d�=���\	��Aa>�Nj��m�*.>�N�+�H
�'|#�r=�IA-X�g*R<>��'�zl�����X-����0򤰹��@�?�r�b?C]�`&]�<�{c��d݂�E<����D}��Ut�l�P����Ơ�?(�K¼DL�T���Z_�����`5���]��a~Q41���)����Q�~d��'��Ϊ��Ni�R:E��f�������>J���h<�4#�~����à�uA��ۜ#����^��3�F�k������^�`"�ѹx�ٰ9	����?�=����@��"��p$�zB^��mM��UHL���˅<��2�%n '�) �PիϡW�[�S��i裻��!�a�/��f+�n��nʤ��L���_w���r�v~�ha�%3R���
�=��a[�]����2 ���ْL��q��CUueeQ��PJQ�ڪ ���nL�"������j��t���p�	ǒ�h���)�OƘU+Z3#y�`0��%GA��T=�ח����.8���ǡ��ܛM�o��#��!
m�w!f#kD��
!k6.�DFA�0���z<aj
zq|�I?��'T�]l�&���0�/����:��K�S����bJ���v9�/�ԏ>V% ���E�y�����!lP��pߍ��J��>U��@����I��<����phܸ�8�.���� #`��U�%O�;����O��o�q6�Y*����`(*��K\�zg-w�b�OZ��$B|w�9!)
Pu�����KQ��E�V��<hd�f�:M>u@�����A�j�=��?�P������%r����؀��8
�Zv�8��-�Ϲ���HL�Q�������F�L���b��
�����[^nj��/�Z�)LCI�B�@<zc���L8ؔ��������q^ ��{B'�~�{�h�B���"��]�ƹ����3��넣5C��41?�#����G���W�K��F�\���qR�xK����6e��~��@b! �CS�h��,p��o �|�,�R��H��vd�Y`�#�S�#�A21^9�eq8���O���t��	Ԁ������
(�@�g�+�^qOD��҂C�`8����]�J�JIU����7���er�� �}����Y�xN��cC�ܣ>ƫQ�jdߪ8na�B�j�WzAS�'�=�e���Y,9��t�?EM2��d	��_"��b��J�Q*��ՒMP�(TOj�A�]shg(�:�=���}����s�D�����W��m�t�8�6p�d��S4=.�9U���u%����~���2��"UP�u6�n��.B:��M�^j��3ĳ� .$��?���)po���� �$:u=A����SC���T}k�-t�)ѥ�%n@)�6ۅ-��	�b�P�(�����Pj]lG�$��w���h/�ڎ�/M�,L$��ɔ${���"��6��s���`B@rdƁ�~\���x[%|��K}S��te�ɟ�)iG������8c���SgP��F�a��2&�>��Ӳz�H�ӕB����P{O_�g��E�	��Ap/1y�O�س�)[�[�)� Xq(�[�z�ME��5���Qā���X���Œ���f/�e�^fs^�ު�Y`��p�:+zT���>�7�
��Z�dr#&��bd�ǯ�$:��?��[��2ݘ��,��mS[������g>�]�b۶�s�H��Zg���+��ȴ��Kl�������m5��1�P��t1{� U)���F�2�%	��-��/Gr;��8A �FUF$�ՃvfV�n����+^�?!�o��<z�1qз�=K��Y�5���RTek�
��kUN,��-�s�����E/i�
��b�ǲ긄W�1Ǭ��BPJÚ����߬��uN-��<�i��Y��+�nO1�����!�~��q+��^��}�S:,�l鳕E6�[c�qH���ѯ>����o��1_�S��r���� z<,WU,��z쵝��g�@��c4CHp�Z�Z�4>�ۙ_�\U3+��0 �UV��I?�衛R��R��v����<M�7ѱD֣���y�e���wguG��M���
Xi��\���/���5^P�)U(]�o2�=`�tsO�����E��ô1�L���=�0����[��(F�]��8��:V���A�h���Y�"�m��{^�D�*<�&��`�+z�TF�p�H���U��^���r`C�@p��.ǯ��h�WCF��8pR�'�덬�?��/�!�����q�f:J"gPF�mz��>��LS��58|^E\��u<�Y�2?lL�����UGs��[�Ysqݯ�P&��&c���e�9�]-�����Od�'�@>�{I�H����4bR��dMԒ�F��ӛ�Gvن�Dyn ��/[�Q-�9qGٮ����u���v2oj�\���#�=w��~�>��?�ҝ���!���^���yo��·�y%�����WYݘ~�9e�(T�3���
���"�"�eK�oI%X��/�V("m�Si�ˉ�F��� aۨ�;�l���16�gt������b$��No�����`���B�C�]A��p�ut2G���m��!�����:�Cr��ti�S���$ɛ+:)/D�x�,C���Ȉ�J�.�D�_��F�<o��{�W���H��C��~鴾���R}���h<ɨ��E�d�g-��ު�-D��MYj��,�d�Y��Rٯ��wX��f��>�Z�`�ҩnS�:���]P!��`o���L��V��s������f�"��������ε��a�s�(�~dr����$�^�V�i�#�U;�CC����En^�S?���9�Ţ\��B�D4=jW_V���9Gh� �&(�~d���.t���	|�{��e�ä�4����fH7�\W.U��R��]�8��N�!��K�����B�	M�R�d�����US0U۩"^�5�>��K��)!�?)
��.!��!����.�/���ݛ�/2�T)c���{��
E;6]�O��Oi�3[�mV��R���R���"��L�BS�p$�F�Ja8,&4�	����X�H!��j+e#׿�(�%�桭�n�߼��(��Krf�Z��C��Ꮸ�g����|��ʧ8
fp�?WSr�ȥ��g�>9�I{����ͧA�Ċ[%iL/:��+�MC������2��W����ˏ��Mg��R,h��I��Z\^�D��2A��Yeu!f:%�1�Ʒ�F�z������)=FP=�ʚ�K��絷0o�N:�#����T�sE*�L=n�����r�H �����6̀1��@���hM��E���4V�ئ���[Q�nH��0}��[*5��C�`{n�A��Ђ�w�/�)�kUi6G���v&�FT�(�r��`-�~6ReԢ��+gQ�Yߵ�ل����X�j�-W����'N%ܷ��̿O1X��"$S�����pjX�1����@3_3�*:�f�7�΁c�u7�ˊ���u����b쏜L��Gַ����4���c�I���\���g����"K2#A�_�񋍪��4�k?���\�/V\bp�-�6_]N�dT�.�ӧʺ�ҝ�*��c�,\!���;��j��bX�D���7�����5U�iP�@|r�
��K7K��,����ģ.�n-��
��]��J��r���S=���gR��8Q�S]6�ӆ�[|�_E���l���W�H&w'�k7���F㖰,������L��(Ɵ�V��
�]�-�ɮ�u��k[����Piؾ���)kf�u�H �M8?ٻ`"�ɾ�[@���O�7��|,���)� ���{���6����&(���"b�[n���>��E���$�:�\U��)��16UYA�^�d����h�/O5�����
	A��>�O��08���W:+z3v�})U�q��$��H��RC��'B���t<�9!��nn�I�io��lN��y5��d*'����j(_�Xd�a|~6:�����>}�9(&M�I�"�m�hyB?�~0d��w�\��Š����H�r��������0Us��DBgRYQ��(	�!AF2�`h�#_���IQ"'yl;U�^�K����q���q��$8);͚�cd7����Q!�D�2����,����ln�Q;ϤXش�J�Ӂ�*mIIc���.��z�G^T卹Y��m ��;�aB䳌<x�q�E��^�Ցs��,���Ð�N09#�9<�_i��6�F��f�"���My�!��C�ۣ[��P��m@���_$�W���[U_�gC顈�B͓S>���
�B�̼𛩭j&�=V�n��LS�dl��ҝ��?uI�&~��*S4�������l���!�ޘ�q�_�/�F�@�k�F\�C�8+������udf�DXU^rÐ���Ry��0$$q��z�݁��К#Ih�o�	]�[��m���Ӌ=�M�&ě�xI�c5�j��d�8�R�
y���qD[��)�gO���t�Ok���ܬ��g5�"&p��
z�,��W�uڲ[[�k6��,��P՝�'S=���� sz$�h���t�!z�k�w`����r)e�F��?�O��u(�	6eT�Z����-�:�&r��(���@F7dyO^Ro�<2�BĄ�j��gV[ۇJ
��x���!�G'iz �����XAN��k��Ә��D��
��b+���·�1V_�H�����KB�Z$�\J��\_�m�����J�qhj�	B������ڧ�E�"��ĖB�x�''v��(�O�N�[�@��
�I�Rڑ����N�Ф�Q?u%"雉��줦�Z�w��;��@I�U$#P�0��w�#�3f�e� T�&Z��v���1Z��${��H����gk�o/���O<��;����f�m�@���]cϋ��ԮSdn�M,۳���BKP&�M�'���5?�s~r�匜fУ����R�Kk<C�#��h%T�@�J�o�k}�CT
�ߑ4�gK�,+8j�
t���.�t�U�,��I�F�7���#�̈́ O�~�=҂�Xs�AT�T;?���W@L:��u�e�0�g��<d�rB|��2p_�ai�x�	m�m����B,y�0� e�IR.����#����Ӎ�HU�n��[�G��Gَ{ꉈ�_�N��[�Ԣ��5!�V"7�.4���o�߀QF7"��J�YC̂o�yB�� ��gIi��6|����4'�NU�,��p�y�S���2L�&�x��m9��P����	.����s`cȚW�����Y#�r��)N7���g��M�:<��Kω����mc� �����]��������C ��j��|��T���<:g�%
$��[K�O�	6?�`�Z��j�5Q�8��a-O�އ�$Ѭs�
��Ī�wo�+��D7S!W�(L��0����T�A�#�Pu67�r��gz���L�h6?���]�>_��Z2�d��˶7&{� :t��&o��V�q�_�R|t����'n�c��0�Ɩ�AI�:hM����~x��ξ\��ͣ":��x�*��)�O���P֚<s;&Vm)3�Q0#o(>���/�����u��z��C�X��UD��ؑ��.���B���1��n{�<�GZ,��/z��~�앲-v���n-����m>�F.���A�-�֫]񻱄l*O -D�z�[�m������4�Q�q#���q"ҷ��{o�95n�w�K=|��ٗJ[�D���UC��Q�YB$k(��$�-,����	8RB�ւ�h�h-�� ;��ö?�f�	GM��t�d��>M9�Av��"�Fc�)�}@z Ol��&�pfo�v�0{Ib=����%���:!�HA�� �ja�ᵍ�tl�n�p���t5ގ�jv@	�Ǿ�9��\r��Fâ����Wt�.��35O6dPpp��e�����]�9�]Yi9�a�8����9�����o$�J��x�]�'|�s�i($Z�Uɮ���q�:F7�$jQ��|�L]�Dz�����~�*��ql�z��>����x����<Ŗ�Ţ/ڋ��򴛈����Z�L��k�ghi\�l�'1�4�ԟ[��)����?�C�-����t�s�1)W`�S}����H��@�	���M�L޽������O�����^���4�R�%:�yps+������G��I��N��p�a���� e�s.�&�ǫ9�J���%?B��ɲ�gxmѩ(Kj�ssLy�[�i=��$\Ƚ.��n�c�r����jZ���jB���D9G�����%�TNlAp�Ѳ��36 ��GVGet��X��eq��}ԕ�I>��u������V�[i�	���ٔ�
�8Tv�=(�e�Td��C��P �jZ��0I!�q� .��ɖɮ�kU���Ř��֟j��2y��S�6.�S���"=�����eN�٘X�|ŕY�|a�"ɻá��ɨ�(��A =�a�ŷ��6�w�ی\�Ms�[>�0.������ {����"���y�d��r�?Pyd�zI��8E���/��'�W�~S�.�ih%�/�bY2�9��pӣ����ܸe�h��a��mue\��|~6�Z�4� ¿���q ̀���pwkgS:/�����]A��]��l�R�idUZ�)]��т׮�.�ghك�%ty��Gi�ȸs�0�+U�<i������@M���U�ě���qw7d0��'��}�Q6���
��`�'�)��u�
���?�F���QB�A�L�^�,�&fc�l���-j���xiV�S��eP@��N)��QAݖ�=AX���C���g�5��M`���\Q�un����z��p�|��Hh�0�\���̖���wH_꥘l@3���iiB��J�L��2�/X����JH��OJ�rRP��������ж��)f}դ�n�xU�@�L)�I�0>�h�M۳52Y��Liel���)�$p�	8
ֲ�͘���^m^i` �*f}^�a�G�X�5�C{��PN%�ڥ�8Q|����x�E%1���