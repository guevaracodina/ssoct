��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ��p"���C��T�fX��k�+��)��6�'�3��$���)��2�+�
�#�7��Ib����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0�6�`d�&n�\JNm�țݲ�;t\�7.�4tU�%J�bdR�yԩ)J�-+����*,�W�h|�����8=�K�������7.�k��X}[uZ���)'��q0�1?,R�i��)�,�Pqi�l(���y�'� ��e>1�5�,��&�%y?�1?�D���}��=m�s�,�6�1����;��Z1X=�b���'�*1/�U�����[�p
�v���j�W����@�xP���s>��Q"O�/ SO!If;�&�A�g׍aw���+���B/��TC6.���M����J���6XB/#�����|��_�*�_i�s�!���G����C"��d:k���QO]��N+DIk�_�AlZA��m��ө����ٱx!j�r��09�jނ`M�4SFAع`��)H�R�������� B�Å6�j��룃͡��/=�_�=8��z��*�P���$��H𲫋�
���]^�`80VC�=����E�k��o�oq]�h�M=�Tp�h4�ӈ�,�u�d�aӹ�zJi'Q�h+�;�(,�"Ļ2�j�ڌ�v�63.�����r9}ҧ��x�4���彌�j�b�����������]\�X���OܗQ<��)�/E�A�ʥ�nY�Q�T�D��w�n��'��G��7�iT,����yΌ�a�?�,\V�1V���*��|� R�y����Hǉ��H�W�Z�.�\��.��<01X� ӆC9�C�U� �ҿo�c�Sڼ���AeN����W�K��mG�U�MbF��;{���M�����pxGR�,�2���bc�aSU�m*�a��L�; d�[��!�62�:��<�Ԟ{�x��I���4Z���fC�"�7YD��u}ۛ�5c~5����wT��̲�/)Y;�������HWԤ��_^�K]�ڊ&�p}��/.�q��Q�lII���q���Wb�2�D��x�bx��J ��������? ���35)�j�ܐ]Xſ�t��[���
�� �wO��>��1�찘���R�NXW'�t��;\X���̹�P�u�/�'�Σo��bP
��cbe�Z�jqT�һ��)X�v�K��Q��t��'6^��Q�&a-��P���*)��-����rf"�g
&����
AE�-:���;��sȪ�lͼ�:`|ەT����i|93������jwUV���w�`��G��ј/G�PT�fӟ|XD���fթ���y��}������s�<r-7}ݨ��PH�d���ݎ1����x��W����;yW4���=�z�br{��u���qq;��Ռ�רL� }�6��ӕ�MvÖ��!��{)E�v��z3#�K�]��ga{���7O��
:٩�Q<��=�`�O�4��^6�稯h���j��d�b�� ����R� �j/Ȅ|cJ�'!*ţ���_0D�(��̼dV,�O��űJ�FL�[���/�m�;|�;�i�!� Z@�_�2�S���;��@*�u4�c�h���3A�������,{>}�z�Y��av3B$�#�`%�43i������>hI.a�o�L��̴]Y����k�n�|\�جj{F���x͙�8t�r��a�M��	�����Ȁw|9�&�$�-�H�[�*7�6�|�,>yU�_���g��� ���-���CcM����\"��e������O��Т�U.]~�铏~@�A�G�f�ŏ��s��~�-�e셞~8�u�Ǭ#��޵��e��f[�pS<�V�je�, ��R"�e����x��>��E��nWK"׾Žn[�_�C���m�-� ���v�AY�ٛAl�6�ҵ�w��\�%I�nCn4���$��;���j<�K�Ρۓ�}����^���`6%uԒ$����AI^��Cp�7E��!�\H���yB��X�W��jj@�wn���M#��b]X�8HАm���FO��6���L���_JF+yuM�>'��0�#�\���7����F���If��'
�z�ՙ}Z�T*�r�^-i2[����u�^ |���"Wxs�دf�pȸsOe� E����\�U������W�a�t|�d\��D4
�mR���{�l*��X�:,�BZ�^��k���1z���\Kv��@h��!��P��W���Z��(���͡����<B��^?˔m�}����pK�f�NB;�`|ݴ�b�t�lY��d<�N��܈��`�W.�"V˙��Q�u,��IY,G�ofK����|���F''��19��R@:9�u�s?�Ԗan�[�8揠m~4��A�N��ct2Ga!M1\͚�m`	��*���5�-����������W���A�o����u��֠�i�"ĩ�5���J4^-��v�,��&zs�>���w9z� Cz�s�+p)��|55��8 PZ�޹b@�n9�P�6k:w?�
8rF��v����an�G���'��;YȪ���y7�:��&�cV�*��(���Z`��F){�{�ڬ�7?Jl KJ��/�d�v$���|:���e&��D�Lܙ���Uʊm�����	iX�'�l2��^���@�mL����l�=m"����l3�d�2>_�br����rU)�0�{[ޠ�}z����H	$L��ۄ�$�H]�����
������l�TkR�����>�.��	ea�g�
ڲJ�癟Ƥ}�R�{�1#o_�݇�qf���47�����*O��kT"�T����wuP׭�GW�!S�ٍ�⎈����r�%�i��Z��U���S�45�����ε�\�d���'�t�9ډa���L�����!~�=v"���7$= 5�E-����\C*�O[����hb�U����d-A��G�@4�ͼ�j���5E�o�E�}ѥ��)���KVF�$_�f�A� �+Z�L����V�+�<�����0|�����U�_㈤��a��6s���mn ���_׀HA�4��ޤ�7y�@�TC��q.[��V���_��lo����Gk��������ɛ��`ͫy�'t9��ӺL�u����g���՟��m7�r'��D�m��7�I�@4�$?&PYA�(�k��?�5x!�1��� _�����x\��i��̑��l|%�8�-�I�^k�ݓ�դ� �ج[�C葩�jઓ�V ��n�T~�e~Q�}A-,u���	�Ǧayɿ�nZ6>rD{�z���w�
U�` 䘦��k�"'Qȝ�6Z��1}@am�C�S�]"c�tNp��Cb�,抎{0��iO�R���$��[��� ���6JZdu�4r�'X&T��*�I4�b"�ڛ�%v�g�|��k�k���!��d�1MC�لc7���;ZU�"B9CS�ƟY0��@����
&�_��P�Ӯ�IХ{�eN��=����,����I�UW�W��z1��XT�� O���m�or�L�NF���hH\�R�/^��r��s��͇6�21��=�Q�nG.!pi?�K�+�S�q�*Z.�0��&�<�K�]7�a�g̉�{s�)LN�H�� ]4P�ˌ޲C��N��;�x���=5.1ԍ���g� ,Z�d���Y�7�a��O3��e�h��)��؍��)o��=7T�p4�66�ǡ"�n>^K�����;��7���ݏ��� t�kD-)�0>[= �<��=�OO��><	��H�Av�G��W���$5��<��f&�n��j�k=:Yԉ�_��ue)}���9���Pu*%�%��	�L����
?�bDpZo�ٮ|�8"&��vx�}ԑ'�^R��Y���W����*�Bיb�5jA{ZBp���O�&���i&���䉸\�/����Z!���bޙ������Ϸ�-=W�K2�Ǩa:ۍK����X�_����;���ْ"/-6 �����F��^�:ǶLh]T�L���Ā����O���yO�=���@`��f��m]Fn6`1e�r�{�5�=�z!�cu��\�p`vic��]�7K�p)fX>�pݕ��됺�' Eʔ=60^��?���=�؃�d��¸�������S�a�iFt�n)0;��vn��%v��hҙ�2�*�ٝ������zغ|�o#�L�N|#ȊQ9[���S�A�^'�hP��l$�e2��A�e媥��-^�Lɏ��m�yG�m\X2��{����"��O'dSDM��\=֣�	�_4��6�����Y�E��i�U��
)�w��sJ���.��u�5��xJɔ#�i�|6�u]jb3�}�)gj�4b��`^��r��r
� �<X��6TT4!�Br�M�&	�䳻A���������>Sc�[��}��ϰH�U�I$#�GKpy����f�v��J�1!�)��w!�K ܼ���Y�o�܁��c࢜),g0)0LSR�9�J
c$�ϼ5�	�p+�~�r6צ�����ںV:C)���M�뻋��W|�6�v((���n0�zax�1m�S���q�V ���C�˧1��Gh�;�t��9�|L�L�����%���9y;I�+����L���$��K�AX�I �p��s^'fƭ�YDۏ��������� đ'���f<��C>��=0C�]��
�
Xf���J��M��c��J%_��(]�ܨ�u�I�������U�#�i$怑t�K9�Z�j�֒�Zo�ou&��hK��uu�D.�rP��3)ɀ �W�q��z�C�T�'{F���2)E[+��*�3�6ޠh���BZ���~����۝�f�4�0eֳ�Muָhd�ve�K3Ϸ�)f�K���FwDrx8� ��q�߻��䐀���lu�C[��}*حT�'R���kvÄ�3�
e��+�Q�F�fM2$w���~Z�@�֤�K�e}B��^��1��?�j�Od����4�0��2���T�6c��0�.pQ��R�#�?��Y_����V}h=s@��nN�� �BԞ/�e'�!��+��B�RD܊V�*V�)�l<,����l����LFy�\�M<|�Bȟ&&ܽF��$h�B�gV*�jB�gfƂ6��]χ�Ď�Lln,3w0AU��ya(_��e7+�;���V�D��HlR�T���1_�G�&A��Z�R�w�)ɘ	7�w/�Q,$�z����%�M��W%���w�ls_���<L�T�a��MLy[bMrJ���Z�RVO�kF��q��Au�Zu
���������r4Nq��dB7�U;<��$�X�N'�Xc�Q��l��W�gVE"N��K�)��7.��-����:�/���?Α�K�U�2S;D����v�!#dN>��r������M9�."aVH8�\���O¿��	ȦdjzH�)��8OAk�����W+v�/i�>w^ܛ�i=�9�cȑ�ay8�B��|�9��R�l��L&W�1<;EK���R�
��y�#��*m|��+
{F9Z�ۦ�����r#��T���6�����6�S��U��N�X�25��z��_�s^�J�7����9� ��Xj����a�8��-��]�
�m�ݬ�=s�7�L���Ă��R\�;zх78�-w�����n��1A��Tǵ�+�#/^�����W�@�?eL+֙�k45_�\v̡���K���'U ںsm��-���g{���X����],0wݽ�<�� �$5����ty#:�t��1q��w�p��;�8,*+�}W�|_���S��a*.J�AT��Ur�A�̌؆�&�����kI�q`�.�iԀ��?�\>�x�� X�A�dq�)��r^�+��k残Ky�1n�h�s8�"$z�P>�I��)���;��T���4�}��U������zN�=(���N�(,#A�g��ɂ�F#G̦X2�6�y�1r�?�e��E�A�[n���>x�1���ȈfSs�W?q����"����ءCz)�]YG?f�4�_��d?S�����.�.��as�� ���"��s�-:?!� 4��5DZSªE�d����E�FJz��M�>Q�P�r�K@"��v��3|б+������O�J�ݦ�lS£�N����7��|]��_��Y�Tz�~�z���S)X
_YA�+���B7d`�j^I�%�u-���̒J��Aҵ\q&�����m�hՏ��|�'�y�E^7-����(q��J�epd�2�Z��0��R����f`����pR��r��