��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ��p"���C��T�fX��k�+��)��6�'�3��$���)��2�+�
�#�7��Ib����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	������*;���X|`Z�J����$2���C��� 1N�p�;S��S�Jz��UqV�l�Et�S~W��zI�n8@�},b^	��� �7�懨j�!]0��X�O�^=��zɫ+�����!Q��Fx���E�=A���׻�n�ٛ]��?H����ⱅ+����&��|]8��ÍI_��q�������9v��S���Nv0����нR���ft��<�n_���;��p#iW/�^a�@��|Y?��>�G��6U����>����s�a�G�Θ���"�t,1��h�˦wW���&G}�������k<2 ۔�쥑B�� ���&�8)v�PH��ۊ�0s��$�'	���q��6�;C�h��t�����&�xj�\��,�������mE��(1��Ge���C�A�eȋG.�W="rYA��+�ڦZ�a+��$�!��OcE���<7�[���wS�~�q+������Xw�OU^�	�ȼB;�����4aB�+���xzӼ�z�@��1�5�H�͔��`.0i�ĢyPیK�,�'�ç�33���h�䷵)���m�* � A�d�A���7@�Nٱp�v#�#溧J��1�O �M�'��7Qk�}[@s��䞕cm��V/ā�IZ.eX��F|�/��[�?\��H���ԥ|/Z����Y�+irW̩P��y^h�R0��;�yK�~f��Øi*�O�i%���dfľȼ�W�l���n̾�X�9!J¢�}N�J	��KU:D�ig~�S��ڎF������'^�/O���P�_��9��%�m�2��uʑ_��.�N��ؾ��x�K^(N�$��R�l8��4��Ca���`�4�R=2�-������$F~��iU�0��}�p�M((ef�P�j&[$b%8�a@��3���D�FOk1�]�*σ_9/�x�u�ҵw�#W�+B��]��I��f���2�5�����s�Ƃ�9��C�`�8��C`��08[XsӚp���$h֌��q����[j��(c>/�.z��=�"0���E��x�.k@���\��gn�p-cV�IL<(p���`p@�ՠ�0O�4�6G�l���c'��2���4�m�u���5D�L���bD5���9fk�'c�@� ��p/�g�u�aC��/�`(�D�U�PV�T
��tyI��S)Bϋ�@*�h�jcΛF�|��wƜ�W��\�})H�2"�ƠJ�V���9�δ�Lf���~'�Dvj�U1(4K�����D��ʾ�5�b�f򼏯�/��4ng�Y���v�Q�S�qA��'qv ��O`d*�����g�i(7�w�Fa�RYim����5�t����-P3$I�y����<.���B�7J*�fi�@�g�k6g���b»����ט��vC)�Yq�Ts�#J컐> P�1w�/%�[H�C�j�B�Gb�r��/Ʃ"Ƅ����2�1�͜,ػ1�E���ԡ?{���t���Y�4�;޵P����<�ŗ��-8g�l�v�S�^�K� �4�8
Ҷp8h�з��cE'��|`�����X
f�K�	2��fEK�LQ�/ך�~��u%u��"Xh�c|�#��?A��]ڋfKd�B?�إ�&*�	Ǖb�:������jbψ��.�+��s���j޽�PЮ~�Q��'*i�,�!n�����#�����<l#���Z�󠢥��c���8�D��z_�&��+m��NIy�4��Vi�)�v_���hcRJ��b�g���pO�l�W���O�t��� �2@��+a��3,����i;)��(P���ԥͨ�G2G���drz������>|��H��Gś�Y�dpb��+�\G��}O��WX�5��t""L�o�zhf.,��_r���#j��g�2]Kq���6�W`��$�^�V޲`����.!��,SKxO�cP3\�1IȅZ\!������l��$��w�5֝�e��8��A���i���F-�b�q�K��p ��`�ެWj��� Eiq%��\A2����=�m���q�$W,�n"�jp2�Dns~��5b��h]cpJ�x�� ;���K=t�-��Z>v��d�7,��$$F��١����0T�q�7dXz�I��.�Έ�ؠ^1����#˃�ٗ^���/��6�-���̦Q�6!���|{k�	ҏ��6/���*o��y�)}\b�1���Q��j�V���=�U�ф4iph�9�y Іĩ8�'��S���XQ�d�d�w_(�}��������7�r�K/q��O�����B9�P����i�0$PdQ�j�r'*���U�߆ՈB��o���d�0H�oNR����7��1�IZ
����F��j8'���2��q���s+�ȣi|	!���B���M��Q����2}�^O	ਹ,����pY�C��7$�n���+��U�cݾ�:�M�[�~D5��k��:�nz;����f��7�I
h�8jF��}:��x�G�-�V4�x�N���ߐ��"\�K�@���M8��8�0s�. �g`�E�G5Ҽ��	˅ ���A�IuG4p['�#�]��x���ك�� ������c��xN}ƶ����q�+�7��^�%��8�+,�:Y�M���v�.���rCC;����� �Uu�4Z�I����Z� 2��������Hx����$���r$����u'���*\^���U�=l K����Yg��R�����#r㠷��즯"�g~(k���Ԯ�MT���%e˼)S	+�tI{ ��+T	i�C��Ӱ珸�u�.F������D�S�1V�&bl���H�� �J
��!��������o�d�ޮ���J$�� �b���1��mOk�Z���N�o��%/D���Vv+m�\��]c��/V\�%�HĚ�lî�cԇ#���,mkv�g4�<��x��Dibl����)���,�+f�8��
�v���4���������Xa�b-�8$����5)�b��8Wxˎ�H{")�վV�������`9���P�.z��4��~�<���.~���	��]
{���f��8!�k�d
iI�-#aP*��U�/�r�
�b.�X��)����&��!"q���	rMA7j?���	D�W2�_�宖6�LO�Z�f��G���D��@M�'�n�����`8����4�u��s�/�|�[w���6�b�%<2&)�8��;d�9�KQO�+w9�zb�P?�N�}��&XXS]2�����T(�ÌTf�����i��#s�Β��l�ϥ��^D{Ѩ1U�U��IՋC�fm�20�U�Ѝ/u��G��q��@��`\̥Nǆ���ٯ	�&��1W+���}��:ndZ߼D�o�8�B��JJt���|,�jm(�p�S�yYY?�^��
_���sH���c�Υ���ć:�A\y��?.��H�l��%��t�z�s�4ԀV��8h��lRn�(�_�VnN�I�94�+^W��F5�I�8�G}���BԪ�����f������%�@���~z�O���ɳ�q�q����}9]�ܥ��aZ�v2���2�ӵZ��_9�-*b�#�M0(����@�]^CS[[��EE<��sR��Nh.��~t��r:�X@^��y�LX�0=�@�"�Jf�lBT֍݄I���#��n��m0g},�>���'EB��~36���N���}%�#���Qj�'!IT��*�f��*� K������w��aV������;(���V�~3G�GRMT��(�F�f��j*�������XЎ��?�]�4Jq9Q��z9c4��!|F�?�Z昱t����w�"?K����fҧ�3؇�)� ���C�
�@�y��Ya��kn�^V�K�-%ٜ�=��'o@B�f?r��{��¼�
u{�M��Tܠ��T�sK#����N�����!���r��.+�R�{����Wu�D�N4�b�nz�;�M�Q^(z�nA*d�@7x���J�R��N<��/�BO�����r,�9�	I����˧+��t��m��,�8��g��lo��x���cP��5{l��^27�����a����n6Fm�=��2������wy���Psѡ2H���X^e5�֯��
�-�B�^���[C��&/�e����CyEd����ܚ?m^���?������m�f�����Wws��e�(ثH��G��J�b*��n�l��$���q�(��\�:�d#Ҳ���$�x��6lj�BQ s����9��:u���1u�G� �C$��z�� c�19�tLC�S׸����c�3n1*Cb_�;i��r71}��i�V`���k�
Ɨ��K��o��]�B�@ZŦ����|O�Ӓ���╃K�1%P�^�T"�Ag7о(=��+�5t�R�nyp�]���C⫦ps�(M9:�Y~���|A���#��'SZ�W��p9�rmjh��D?�ZA��IG<Z<�4��4$82��2k�{��Nř3� M��vzPc�'��ٳp"D�۫S�"Xnv�2�l��V��^T�����ʷ�(�F�ebN���;��u'~:�a�2	�rEJ�+r��ǩ��0���;6���/�L��j���X{����N諚F�9쪖�W�����'�QK�ټ�eU�T�4��v5n�O�b�H����1��Z}�Q��ؕ��h�#A��1�˷����5ȂM2��p
��5�Z�;�qr�Iv��!��۩Y�'��W՝�-�cYq�(=�Ul��<���"����..lT�P��4�1@��+çԡ%�+DX^�x�*��G��k8w������3���9/K��+�Tq
 ���ɒ&i�AFh\�!��ܖg��խ��2��@�@���wE�q��Y�W_Àx�O7$I�#?�͙s,C 3���rè�ak�o��A[�ҪH癑N�l)�|��le���d�P%κ�u�8���+5�[�p��'\��25��
ݮs���z��f�<�H���i�3͋�^�DU<�P,�f��*e��r�]tLcl��W���;�Ű0�ewqhG�}�?�y�G��,g��+����d����8j��QZOm��L���'أ��^��z�.U�����]I6���:��&N��U<�z3/�5�ݻFOH�P����ho�tuuR�@�M1�}"&�Y�p!% ���lqٿ�-��2|C!�b�ʼ��#L/9�1�̶�vI�kaY��AjYc��ڲ�'�*�2`U3���,8T�-��	�$���V��|�I��!Py߰[�	 hIm�\�E�]�p�؋����-ݔ��u4�?Z�p�A��yΕ݋�۾�V�!֐��_ZZ�,�e�(�M\ 4|�%k�V��$*������0 4�i��P3�l���r��y2k<W�����"Jɂ͋����j6ZuJ`u��+��:�5u�;�nL'SD�Ub3ĥQ��6��O%=0�9�T����(�aw�Q,�8�����'�zL����VMd��d$�o�!2*/S�H��X��W�sc���㯈��R7O��]�P�:�Ӆ[VӠq���U�a�qf��m8j���:ou)Aj��p,���	<j���d9�Yo���[��Q�����X��U�CΈKO����Q?(r���W�F�A|��CD�"���2#K�^�̾_��H�*E��8t!���T����iO��8>t9e�;6��w(�����L��3�ʷy?@Zf{S���i�=8�Ȓ�Pqw���6�ƈf��-AY:{Y�mq�[4���>dÊJ2��8�W�lu�M�hc�b��M7fV^-wm<����Os�6��߹��h�_��Me�S;���_���l[�ᡥ�Y�o-�b�0��@���0�̌h�}�<�FzT	��'բY�n�)B9������G����|<��RBE�nh�G����j!Q���Οu��d�C���K���J�Qmq��!��sz:��H�ő4�ETf��Xp͛�#�r�)r�q�J]�łH-U�`_�s71��p� x;�7�hK�(�����:�@݂G	U�>/m� P+���t���t"m��
��`k��y�eS�v��98_k��`�e��h%��~^-j���"ANׯʊ�u��TT����#�,8�`�S82��o����<�:�e�6.��T����p&��+�'�9�� �81G���L��l�b���h����VHZd�06�:�a��?]p֯����-c����S�(pdK��6��bA��?~�%U�)�p�L?+�nQ[�xD��#��-c��w� ȧ��q�Du���n��:2��MԓA����|�Ϲ�����������,)����X"�\�fV�wi{�:��+y�r/a�&5��9��M�a�QB�ώ	!�o\������4N	��5G�����a�M�^]��v���AH�� �s��������C�,�k&cB=�8m0�dA�[�W#�-0�n�P�N��ҧ�Yȫ�u3�����a9癩&���bNb8ˀ�d�#��3�(	���юd�I��6	��楸f>Ⱥ���J�ҍ����t�^B�}���k*?4!�������X#���\�|L0�Q9���t���0���6��^l���b]Q]�����I�G��l͂t��P�C�5%��h��P�7����t��Xc�@t���@z C$����������AoJ��-˅|)5|辬!z��"ݽ��I��.D��/4����<�)���}����7c|zF��N
!IE���@��wWN@i=�]�bC�m��%D�席��<�t-�gԦ�T�)���<���w���qY�1��6�n�"���]�nh���ͻy�O��GX���P-���=�%Ձ#�i�K�pU�4�Rp�+w$�͒�*F3=���7���_���n�6*t������:�A�E�����4��)�����<}0��}c"�[���GG��\_�\�������/ޫt�p��P���BF��;�S����ͨZ�;z��w��6���:Y��
L��"2����٠�S^�Q��h�H��b����u�NZ���M�X:ط�Ѧ<;��[���6����_5!�QQ�q%����&��Y�q;����ȝ�Wy�s��ªU�&�� H?D"�ģ���SV0c���̏�y�%�F�\�ױ��p5υ����_�.&7Tq��e�9^�-KܦJFEJX��,������6�殭5Jq���Q��#�8��v:��=�1�֯2�Z����5��M���q�բ�qlќF���a/9脛��QV�CgCDc
�w��)��[4֯���1�����!h߮�\ډ�C�@2����1��NK!���Jr�l�7#�1�X�%�����.�������X�C8�2|� ��~ѶqJ@����.x���w?!�X*�U��,g�����ˡ}e�W�a��gBs�D��j9�g�Pb��n���y�����_�����bz��3@se�F{|z���3Qb����w_P�Lf�zM%�����rDCݩqÜ��+8~En��� ��E�mIiΨ��z���C��E�@�0�&��δ�񏡟��w3K���@=�l��{�^�9,�h���#�c����+o��.r�V׍�|GDL�4���'*s�f_����F�N��2�#����xx��\Ǒ�و�-_�3Ȳ�R��ݸ!q���]���vY��V��\:qw����ޝ[�/��A�$_�O
M�g���jx���O�g�i�c�����Ô�L���o�����;��2�S�+}����U��8�3��v20����~�K�I�OZ:��J\��isѱ0��<}�,T-_�������ב:�� �g���S�f#�^<vri6A&@� ��P������ht|�V<x~nw\͏;ʃ�H΍���zʩhB��|�K��zQ�V-��g�G���0RϪ�L���/-2�1d0�0��=Z�� ���\@�oTCu�s���g��f�c��]sG��(>/b���h�}M�?��ю�Q�_�t4k��Zp��ǣ�*e��m�g�����aw�{ ���ľ�iW*(q�B8�}x��,�wzhk��A��m�
)K���=�#�����Fp�c�S5��Z���|h�~t��5��v.����5ۘߎ3�_k��j�Ϥs�DGW����b|7SY�2�/�|��<t���$����Qp��N�p��
}O+���k��l~�ˍv�;�ĎGm��|�i��{�5�;�״�`���Xh���p��5���=#��$�.k��Y�kqMZ8���L�FK�^
f��yM���Sƛ����y~�&�9_�d˷#��c� ,�UR���5�<�A��_P�M�t�pd��K	�*�;�W[��.�>���j�(��W��%�Ԥ��
��z�d)p4F0r1ީVU�����My�O�.�=Zۓ�|6G����vŉPM�������N����;�i���~����Q5�6u���RFt��J��63�hUA�X��yU�I�z�E��M����뗭�.~�Oɇ[�4�VE|9�L(�fXH&��|���"�����צ����'���2��l���+Lг?V!o�,lH���B[���wU�O��;��������~��pi���}y�-�e�T��O�h�i�F���**x���.����C����GN���9Jb���7R�ti���z5T,̑�
"Y"��vk�(Zv|�ӳ�	����5q#?�t��I�<�u�F��i�N�A�'��`��h�C�R�z���^,�?UM��_�Kֆ1牺~,�!�Ĉ;Ǟ4�_�r}���7~q/��n;	���p$.ҳf����!�@�Ӵ�ͯ|�����DK��^L����lc���+4����#�9I~8��|!W����H�u�񅽲��f21X�e}�TM+ζf8s�J�@а���e�=2s���yJ?ugx	������[	7��*C'�F����+ڜ$(Nԭ[�R�2��b��}Pdb>e�5�KR`z63��K{�����S��	�?�����S�Ye�7E�KBX�U'��9D?m2G�բ�l0�h9Q��L���m�}���������3=���6ߧ�r��h�aM���~�w�4Բ	Q�Wb�0��+Jc�W�C���+ŴR\y.&s���wĻA$`~�)�Ɩ���u���vT3P� ՠ�.�OS+'� GHQ���|0d����e�t�o���8!��4���s�Ƈ�[ނ�T&��a��%%���97d	��CZ,�kA;�f�;����"����~;]8�B�~�+N��v��	i ��[2�P�RV��S��d�s�E�x�b���O�[0j���d1z磒�m�y%���[���~VSe�� 帽��S����^v�P��v"��:��~����W"�f/��c��Ob�Xϲt���MU�u��J��GI~ϧ�Y�$��F�ou�M��Oi�&I'c��5MҼ�㐡)"�c��-nDX��'���Q�T�(������|�#h&�����_ti*w�/���<��*��"�f9{������Voe��!��:�?f�Y��+6G��<O����O��7�����b��D_V��=%|��E���)� yt�'���i���K
��8�!�rG��c4M��.m�J��LXǗ)WD�y���xq��[�G~D�4��lM�z���2���J8�������=���K+}Zei�J^Q��qh����4Oz�`�"��L�2��P~�2��s�1w�!#k�D��(��
䘎6������I�SP���<�G���Ά���ݠL�T��f-P<R8�[-���q��R�eCiD�>(���Y�v^����n
��Rc��B�]�L�V)�/ۢ����y�
�ǚ/��E�	.Na �8Ad���r��Qe?�����v2B,�K�t��/(PD
��,-��3�N�zϛ5<�3��/�{��������殼�~�a������-UP��=���xn�eS�ru��k@S�4R�<x*p��q@�(//
,Am�hT�;;�V�&"¿���a����@1al�E)�{��b�Rk:{GP�,�.��G�y!6��'�N!moyK�}��,2?Nk�s�U���!�V�7U�0�.����f{)����������Mh�wI�f�VF��(��TS�����6%H���\�)]��ʤ�o��D���L��lI"Z�6��?�ѕ��[��!	��ĕ��@���eйfD`�C��\џ�*�籧30F".��6hj��I`ݛ^���8��t���Ѭ5��.*hǬht��mp�W`�R����'�(X�/	�Q��/��`�Ѹ�KyIb�ڕc�-� �n$Ӓ����C��\�m4���	���"�K�z�	K5p��	��&;��ƶRC��%2�U��� �S�4�b����:ڬR�w�á֎>��5�Q�`�ثK��W����k^�%��On��\wI�ƣ��:7���S
Ms�l+b��_�'Tt��E�A��Hm���:�Ii�0�o�6" 3�p�F��������mC�D���#���Eo#�(+I铸�ih�bMW����h6�w��&V8���F��w�j�2(�IY������������q��d}�Ga4��l���TS�R����:_`e�2RƐ	��͖"��E�r�80��&���)cD�\M���s�A�Xch�S@Os�ڔ�R��l�j+d���.QB2(tZlmi�?WI�Ŝc!6-�|�H�y�g���-���^/��*a�"�����@�p��ї���׏�<+�3�t��'j��4�3�K��>P�E�(N	�rZ5�3���j���\�AO��ϩ�ąڀjU�� ��0AN��O~�8bصp�N��[d|��x��_#D1��Cb���$2-V���[��c�yV��ǐ���:|�_�-p�v�o�1���ݹ�q�^���v:c#TY�c ߧ����n+I�w4)@b�85ke��}��bV"*b�7|uB����{�q��Qm�		5��M� x���Mr�`�qp�\B�W�M��6;����ޗ��B�w�����0���Mo-�ܭ0���XA}�K��iJ��S0��΂���}	Q*+1n�њY
��|����>N���e�|25X�ɄS+������q����e%�lP���~n�:�X��r�٣Mb��I"����E	'1}���0�b��+��^ng#�߅	;�`R_�[��2�� �;��,�Y���Hv(�BX����,_~)ۻm'���^�����8w=����B�~��RB���GB�ްq3���\m�lX��FyB��/Yo�d��[ ���E�X�B�lX��%n����t�J���� 	Fl;,�E�p."Ԏ*��ېE�Cz\����2h� ��rSD�|�ŧb�(A{A���iP��x�E�aKZ�|��B��� PN�
�G�v�^�󶭻'���X�a�D��/���wͰ�� ��U��#��H�8`����Ϭ�Iv� go��,%���.0Jޔ�x���خ�f���ĺ�O2�ߵ���������Q��Z�	<R��n�C����2-z>&W����U�A�V�IR�/hD�0�\���䲒�)�9�����&�7�_gB��)kG?%��7Yx"ʸu��8���Z�Hi(��X��'��{�d0I��ʢ�M���ا�.|�,��s�kOs��S&���	7t��%b�М`n���Z\�ͼ���3�h}�R�~I9P���Zd] co3�t�J�oǵ��b|�u$�dLΏP .��.٭i���v�Gp�U���4a�v�/GK<��G���=#�?/�؈�e�C���8H��b� ��k0uepA�o��A�5GBq=���v�� �A��inx��R��<`-}ap�������bj�y�)jP��3Q��0�0�␃�(��
����U���i�L��j)@�j�'�@¯�%초���r3��p���8�f��H*�ǒ��6i ج��G��L·���܏��;޷>J�(�+�`�;�3���6�A9@�)�&���;Etii*���[�?�q��a��g��t��t��@������o�
o46K��j�6�䭦�M��Tj�aѰ����]Zf%n�KW������� �2�A�1�4oGnˌ\E�kY)~����X
���6���?���"P�,ϖ�s�ɦ0�.U���IHd�;���d0T���f���氯�]��Y�
m%�g�c��B�]t� �
��o� �Io��[��Q���AN+F���:����`I��)U��p��@��Sտ��l~h.�DȄ�φR��OM�a�m�
�|m:FB!�p ���'ѽH�E�f�E���]����T$e�s�\�����2��Lx@��q�*��/"��n��v�ag&xa,FR��炡P**ٔ�����""��*I�d�3�\7u�}�������cs����mr[Id��A����hn�6�n?�2Y���pJl:����.N_j���I�"�C���ÕFGe����Zgn\����jH��B�'�yܫU?|��ַ��d���#�Ք��ߍD�BoVȑ����=1_��ft�J�I�N�J��'>�<a��\�I`~Pӂ�r���[�.�@x�Ίēx~֟�Pѿ��bͼ���$<��mǳ{���B��m��bc�I�16.)U}���<-�oFP�PQ�:�ϵ��P���ņ���U>{�\�L�y�3i�����Rzd��>�2v�Ļg	6�u��4$��ل�QW��B��0e~A�i��0o4�d��TXtn����g��4hf� �R�P��½-&���^	j��8�b��$y#a�[wj�%�cȢZ;��\�ߞ�;(P��ހ�ºRDq�š��:ꉆ�� a�5,־�0�܄�f /��5�OW�;�F>.5O6��UZFU265Y4~\���Ŝ�;AH�Up����A2E��8#5C>�Bw��?C& ��ӷ~��K��7���/W������-����S�]��O�_bepQTU(2�j^.�»�Q��*�.f�?�B� ��ġHW�NR�e7���K��Zlb���H0Kc�� ��*kF��w����;_��e&�(Kxl�ɻ�Bt(�o���	�Zi}���H������&N�O�4"����{��IYx|A��0��8��Y^@�'�>.Ԃ���˒�S�0���E.�܇gBS��'�to�4�z�.|�c/|J����]煞j���J��p��R��vw�^�siW�f�N����b�n�*iXN;�mkI��nD@X*s��(�LxT��\N7�6���x�<%rH�W�3���+��U���j�LW�l9~8�	؆�v�e�QU�ߑ��a�PϨ͔:��k�m�����$!����AQ­]�8����2�}$���/��2�L�+3���A ��$��A���+��W��N�Y�Q�	M��_���pO��gm�⥤�����]�4�#RJ���Y�8k��g�L�����ӌ�{�_�9I�^�����p��dt�}��3���!py�cO��6jzr�]F�?�r(�E����6�~�a 7����}��T��؆�nl<���1\z��xe�=�f0D��}n���;�\�$�l�O��_c�;x֮���خF/#��VHPH�����
0}{P��7N�$�~8Eъ�e#+�Ш���<7���a�2d�eJ��MY�>���	_�|A�(���i�p7���O_�턂�jRV.�s�p٧���v6����ټj�.'A]��p��c=��~#����p���U).��v''H�eC��Ȭ���|�|ư���Eio6���joS}�IS���� ����:fv�5�#r�(��_�)�>��d�`7�v��]�T�W��σ*��#p��Ѕ7M�z�Ȑc�G��YY�<�b���nS݂D1zV�;�_�Sl��_��`�r�����i�75����;��6�����M��+��K������G�FF7������-ƍ|]����v?:�����R�h�6���x�+� ���>_�I�+Yi�`�r)p�`�n�)U��l$�D�;�ܑ@���xM�}�Y5F*κ/vj�_�\��2~�`a�^�w���Mu�b
�SA���[__��iN�����6Ỏ�jM��^�	����]���X�!�cDe�U����&�}�����z4�$��h|_$	C�[ک�H�!O���չ�d(U�X�����I.���,����J�b�,���
SlqM�8
��]%KOgWJ���KEpP�×�( y��JPn��,3�$����f+(���WD���UM�37d#TV.�;����D8�����F���YE�jfd����M��2l�a\��{�FN���x�^���q�6�4ڷtڊ2n��2R��c��P���g"���gI�Pl��6U]^�wwui<�Z�����O�gj5?):�;_Om����#b��� �n#�L�J�7�D;�$ڴ}�>iNrN!�A�_e�*ͧ�(u~�H8Bp6�l��L����M��d�9>[J��D:_}\:��zo%�9�&��s����s3���T�Q��@i�Za6�(���l���9j�TYBݛa�?�-R�hoI�;ܝ�<{Ef	S�)Iu0�ϻ����lI��g���F��R��BK
�t�_u�|T 'X����-3ɲ�C����?s����Y3u/����?a�G񞖈�(����ǘ�塾#�k��&5/�~��Ҳ������cۏk�����B_��@�u,�n��L�!'TE\8z�������0�򺍺60u�����6 ���y)"ى�D�wei*\�����n�l���d���':8�N.h�x�T�bG��L��f`쓄�v��蓏�~ֵ����v~4�G�������H|��c�b4Ǌ��a����ue��s\����\]�i��>4��-8�kQ�˃ebU��a�p������[�2����u�75��z�p\�?���ޜsۊ��VBs�IT�q�	B��l�+pGowi�- �
>z������v��:��f�Zu�E%Lq-yQR��&�X"��T�8���6�X�tFՉ�1��O9`�V)��]�?���2Tv�`j�`����,7�c5����T� ��I�㨬��a*X�<K
��	٧��@N8m�����*#�S�(�Iba'?�YPɇ��^A�#���~گ\���������Ȝ��%;H��Ƣ1;7�-�������c�`y��h����.!n�������}�<�3�1�$�Y7�U�M�*�������<�׿MV�nP���zQ;��ħu#\�!2#Z	V�CE����q?���w*2վ�~8�^���iG���-e	dD��{�C��k��r	,m-�#˂B��cw;��;�5��<����b؍�Aő[�e+c�@tƷ]�����3l��Ք̕�p���DRU�k�7U�˿n�4TME�e���=x���b6��"=�O��,�`�X�����M�lȇ-IB?մc�xaK����h���L�2�1���[���uz`�!��`ϣ.h^�� �YщӉu��K�HL��*�67��{>�iKzt����ƺ��.���������cQ.�V�I�?8�}�ໟ��c�靦������Ƿ���H�4�,Fp�*&�:�V��&�q�Tko�c��A�RN3Ao�I�x[�k[q"�$��x�Xs+��C�`^[C��6~�'�)�۵K�&��G����u��l{0`��kt2LAײ�M����d����l�n��uW�zM���Y�䞖�_Z�(O�GU��5$g������p#���?���� wY�t����b V�;�8<xL�0�{Ip}
��D4�Ha�� ?���*o�v�����DE������:~��<O���CR �WӠ�����`�Q��`��L�ܷ!'�2���$-��ګ�ƙ�5Ln���;���QAqC�����E��T��+�y['��!vɥpR�/���,�l��1�Eؼ�;OZzc���7�s�q$t�˚�TkP�\�q�#/3�|74s[3r�t�=�v���1���%�I(���������x���i�=R��U�s��=��Bl�V�5%�eA��;}��+�|�O�
�����-l�S�׵%��*�f�"� F��y�\Sd(����%���+7���C�acN9�>?�BV�vO�S,�����XA�GǞ�)�M^�l�1�	O�t�M˞�m�m��SH:D��vz��R�����TI�*��( h��m9�'�+��^g��r�}���D��c_�qI�\F鱘I}����K
�"����[j�����=�S�jl��{o����*����2@8z���^W���y;A�X)3zNl�7��K*�H��W���+���j��P��9X�Û�k��3�W�S���Ҷ�z���+f�i%_��T;��ڪ��H�edڑ�����\+�8o��1��#K{
�-�0f�Q��B���;�=�7����E/	���b���`Ŭ6���/�	tC�_�P��+�A�Z��$[��U�齋�|ڷ������>rъ7ï���<� ��&2D�^ift73��!�!��v�v��C�1�Am�AR��KOJo�����o�����X�_�M�]��W�[�_����ׁCh������N����{aT��)F�a9x����o�<�-I�d������'��Ӈ�j�V+@�4���<(4P�`][���ODQ�u���̗Q�@m)��ږ�r�J���rDOl���Cl��>��A����e�(׻�y[e�E��U8Q�<Z�67Emv1+O�&<�p�US�3�՗mt�ζ�Z�G�*���{�X,����a`m��V0��iM�h_�Irj�VE3�����e���B����[��JJd�P�kt�s��gc�����"uW�b�CӋ�`2�@����8iQ��tAF#�˱��|��9�Z�:�$�h���O@v�e`,��o'���|��)M�7��v����p����$���U�����yF�e��kJ�Ͼ �9'K�a���eغ�k������=�5�܅>)��!Ie�h�a�"�ˠ�+��Ty����~L�	&%`uej�R���hG&R�O��-u�J���7q�6"�ʱd�� �֧D�+C�
��~���p���1Bc\��'L�H�=��5�I�.Q�B֊��9����wY��T���-���L�N�tBd��ɭ"�p�JQᨺ/-��5JX���{��
p�&�Wdߣu�n�`J�,v�F|=�-+�֤�fʎ@�E��ȅ�����	V���H��ªx�8��҂:������,%��F?❧�����6ĸ�PCO�P_>�f84|�ER$��Z��Nʓ�<�a_k"�Ǖlm�����+=�3��t;N�j
��M�Re�޿�/z�������.�g� !�!�~��eq�~�q_����0�觍9�k-��<ϣ'�J�X���U��m�{v-N�%�W�Jd5��3Yz��e��.A��WN� ���"���$>7z"g��̖����dM��t�u�겠���G���a>L�`o��0ՉSP4�#?�KT/K�2����)�K%��jq;<?/aY�C
��m nNKoֹV�����@. 2X�Jg�O�rE)�#�xGq�U70�\,���� @��]d�q򌭞c~g�"H�l�7��{HB0���Z�.��v�saP�*@K`��4f ��[�q��!��Q��OZ���Yj���/�N�U��ͣ��`�oUa{n�������T��an��A�Ve��K?����,W���R���>9������~�0���z��~�~f�F[u��]��?@�u�FO^T����9Tt%-���ծ��� ����-S��W["m&]�S(?�¿�[�N��#��$���t�bU�v�΁l�F���(�˲t�Wd8���s�ݘyԢ#8X>�(,Z+L G� ݎ⸎��ݝ�*3~�_�68~����VQI��1ڡL��q��ӜQhjK]S��������O6ɚ{
�K~��:?r:`V7��+P���1���{<ȋg�Ռ�\��R!�pA��	����Y���	e��_��jR=�-m�Zd��>n37��MÝK�}gԣAd�:�.)�mub5�	���VZ8MΏ7ߡ+�i5|#ݝҳ3wZ�S�N�k��!��܋���M���])"%��˹�7�~��m8V8H��iHß\�Ct�m�d�i�%d��tSz;����2��uˁ�C�;]�t��	�k�P�����|T���!_A�h�l��z�ri�2�Z-�ŏ��F��!Sz��;�6[�*0�_�u=�r�Y�d�����T���}�rZ�Ei����4�?�lK�[,���ߪ�$�z��Ue*K#�\�Ҙ�1A�x�a�����ަR@b�Ќ���ir�.f� t���͋ͺP:g-:G�R'��{"�3	�k���Ԇ�}����Ł�g.�.8K;�E�����*���Z�dݞ�5(����c,lˉx�����-�F�f\TT�cX5d��H�B͟u'3�����g1b��I�s�
���G���CɍjӺb���#j(S0�ez�8d?EX��|����;�E-l��o<z��gV��H۟c��͹5J��"nv�p�K=�����.�M�Ԟè3��?�G7Q�j�L�cLjE
��x3K�f�������H�̝x�M�[��̐4wku���2K/-Ϋ�(3�;{ײ�?JR ���(왛�4v�@���Ϧ���#���<EԂ�5�/nCV���Ѵ�(�P<},몛] �Dv@3nf#���9��B�'s��#����^��7��AyG��3)F�E�ot0��;���ˑ"��^��13i�0F����~��fЈXrh����i��l9�� �Z���SFF�g�rZ�Im廩�fd�w���V�T�h�yoI1�$X������r�ڸ���"�1��\�K�*�JvP8��.*q y"�V��Q�uҴ� ���+���"3h�e���G���)㆘���>-���B��y+�QaY+rHpЌ����ч�i��5k�=���w-Ԓ���3J��!b@�Z;H��I��1sCY�sd��H;pZ=�w�i��BNYՃ���i^����dS��`#��S+G<J��>�\
tl�n��j?�����.V�@B�!^�K9���رB�v,����=9��&?��;c=K� `�!wHfG�~�w��i�����<)Ǽ�I���&�Ѕ��\��k��γ�'O��	A��L���Ua����j��N ��s��a��m�,{��P��< ��Z�TTS��I��wf����]�	�1o��苆�G@.a�d�4�ӒM������|�j�v>�𱉾C��ʵIN_���ߓ���cR������֋�9�S ��L�^�jV�z���q&qcݖ�c�m&s�����y�)���,���:ٍN���U_�8�y��،�mp�{6	#Y7��>X|�
+m�S����	�-�H]/�D]��T���+��<�@��^�) G�k�6'Y��I�0�ko�='q|o'g��,N�:Tw[�/�\�9��y�_��ؑ�J������;�H��������	}�0��F�ٹ��ႎ�/��|����m�|�̂ms �K��R.uPno2��~�"�G`!�����P�_E�`��F�1Sn���*�(�#���2:��:}��1��>��n�.��%����l�b|�0�X�L��q*jb;�\
��ME�>��:QJz��d�W9�Թ�Qp�E�fi��|��� *X7J-�p���t�8�K�4�@9h�f�����;-�![S�g��a�Z2IP�j98���`y�7�]+iS�%M�$@��!�ʕ�	�P��g���U--ߤ5D3l����Y�N(V��m�f "߲����V%0�9)䩣;���f���Ut��Ck����Pm.D�`�OS<�|��0�R;v�j�����������8E�Ń^��4A������9�5�qk�n�����~j&5R���� =@#�̀R���c�i�g�<��� ��(�	)��=�wc$�c�����}�v�==�3�|2�/��p8֨x��z+3�@�$v�7~TO�V�Ʃ�?!x�����uN��*��ū��i�`� ��`�j�D�>LŐ��t��;k�l�=�0"r�*�w^��e�\�S��Z~m��r$�E����.T�"�� ?��RJ���� q���vm$�?�Ɵ�io����(�Y�~z�N����cf2B\u�KO}���Iw��"��jk�_�[�]њ��}�j`�"�N�A"a!��~DG��jr��_���f��*<~9G�g��^�J�(��r�/�){^}<^��,�����|�v���)��K������`1pd-��NE�'�՝�~P������,��W��4n���d/7i@X�3W\��P�Mxx	QF6�2='ԉ���*xN7�n/��fS�o-&����iܫ�v*��
H5��'Íc@��ݦ��`�探x?��Kb��ڦ��&{��K�#B9�>Cb@���-��W�Z��IvE��٘��&�+��X�e�#NzN��?�j��$�W������g�g&/�S���Pi��vf+�;�]����%�? �����+�l����#i�����A�t\%�6���┕�5��XkL����ØPa��Z��+�:�m�S�/��t(��Hz}4(>��1*�G�L����HH_p�vT�4�'�D�^F����e����Ǐ���AO�jf3e����ڎ�xyf����?ɖ�2�����(���i��U	VM�s�6���Y6�WK�7I:\IS��f ̐~K�^(���F�^X�,��4tx`IT���LA"pi�ni_(<OWq�dn�b��FPL-�!����Zn�32�����S�f���P���U"0�x>}��V��l�������]�S��9����b��ICi	w�Vl0�Aٍ�l/m��6�`����CF������͊er��CY/����U�5)�H"L:l�pޅ��Z@�s�x����^�K<�L.i ��f^f�V��GFۖ4�c�:�{���],CI�y�w���k�HU_�eNs���9>,��P=��\1C"v�s J�̏b ��_��ߪ}�ݗ�O��H�L��cWV���;ňa��T����I?AIBF��r�*#+j�k&�����e���A+��o����;aJ#KB`�A��ij�I/v����^�g��4k��2�dE0�B�͑�fz�rB��+D�,K�龝"j��k�6�`ǯ!Y�L����̗I�WJ�3�%�Äy��y���.��a�ѹ	_^l�Չ\���_�;ٴ�RaM�Q3קH^�.Sp�P*�?[>�C�����T��	��\��Oy�2��F�(/�9����&S��/U�eC�w{v$#�v/���3�.����7 +B�m�n>L�=J%}'�i����\j�=B0����:Ż�OHN�2F/c�u��Lm�Y4�F���Q�,(�V��7�{ ���b-aڗ��}]��#�h��ȑN"|��AXƞ8�j�.!�Um��Ĉ,g��C�ZYn�t�!'5�����̮z-9�� ��(��De?Smk�����qc����տ����̶O��Y�xD���Q��j���lӸ����.T�;��?����$M�����0+e�UHO�[�\�m�\/�/m"�� �*�G����V���ߧF�B�Uy������3Yy%
ĸK�Hzrp��z���H��,E�(:�<�q�`D�ዡX;���E���Ɖ�@�%Xx�f�~Vi��?G��
,�iL��]"5����m�d}��i��w��r�S���|����~^9���\2�3#x%���RQ�6x�cA8@Ίm��b#�7 �lj�&�z��1��j�@��E����V	T�"�L>WoW��0�o�g��V/��$�-��0�FTz�y���"q	��Ϝ�C�Q�k��|��Z���ـs/�;)�f<|Fb`�jR�Ec�'Ǌ�(�o|�9�N��nS^[M��G���:M��� 
��bL�H��Yg���ZrME������y�%8����z:P��Az��r�S��m&�~�D����(�h�nK�cz�,8ѣ�+�\���B�P߽�8����8���b@�Y] ��}��I�/�>�2��Pa)xtz�BSi���ע��}�=r����w��ah���6O���eK�T=b�/�+�]���I�;�И��I����\���/��S&�����΋:W,��i����.�X���=6w���FX �Ґ֟)Ey$I����g��an�)�{����i��/{_�t/K~���^¢���iP*�� l�A4$ѓy��A�8�`�C'0��8m���4�D�Dh+��
Ȱ��/,'��R��Ĺmn�toȷ���cm�;�u����ʑN^�5ࣷ�=�qA�؃�!/�Q��GyH����ЯiJ�ܺ�=MH��r�D-��1)�l9"���͗��'��i�D�X��a���@�X�&���0�>cv�3/��D8@����t\��]�k�M���_�
��oNY�ĞV��O	���y۴�+���<���lĚf��~C���0k@'G1Zl�,�XV���S�P�y�)�vE���<n��X��Ø��f�)�X�)m�ԴmJ	*�XX�^+�� ����5�� ��� ����<�R��5u�%�~�A��tNX3s�D��M;ѳ��a��]\�BT?�t�̔�YvlX��=>�ej~�g�*y(�Ɛ�d�	m��{Q=�췕�N��<i�������?��П�.]�Z��ݺc�6�5�i�6=˯
�
ax$����H���pnd�)� ߹]�ʬI�od�V�9��ȴ����g����{�S�C3����$�}jsD�Y�<���縅=^��G��#���"HI�ZV�5������"�w�hFfY�%�~�0#67���6�Nk�/���ǈP�'n���1%Q��"P!i�����{��_*���Q���$t�#b6�ՁV�߷T�\W(|��(���mT���x���((�I	|�O̯;��C�`��/OiG�_��-	�yS2<h����H+��Kh��&j�e�3����8��M]?���a���v���Olh\j��#���V_F;�?��.l�T=�N^M٢�9��p�$�0jd�Ϋ	�^���z�v|
�PF�ۄ��ΉD}�>3�����/@�DN���xR��C�(��$c  ���"���B?c�V��z�u�A�}�L��e=�����]`m��P��H\�u����/.OX����Vê��Ҥ��%9�*�`^��Y��pP���H�9��N?:��l��>�<����N�mg>�����꽸�=���E�Wg/� �ݷ�S�P1�?90@XS���-�Z�i9iFX���+�����5DD7�js��rf�		��,2������48��v@XK���x�A�Pnh��_�O�4s�D�5��*���)�t�~�B1j�E�tR,�ei�#t�����­�:��eI�n�U��ҫ8pI|#��9S#̶�P��l�&uM�2N�/�z��l!B9$S���:�"���ﰬC1_�M��>�-�H��� kIG����ږ�+�+6�@���Gm�ϵ~��*���N9��`ߖ2N����l	5̔�h0�|#�����	RZ)P�N������`��u_�#��I�Xuk�Z�= [���O�0����p�[m �c���6�:�b��|M5�|Orp��K�e�`��&Ѹ@�ˌ�`����ڭ�Jͽ��=ĳ�e5���+�Y���\��g �<��*����^r�-����b���ٝB3_�1s�`7�dP�6ަ�:YP	�ͻ�E��7
�Tȕk9�|��
���YsL����bK������iw7������D��b�n[�31\�z��������vOH������!�{�{�*��T�`Em�P�~�I�sP[75x�/�}��&?+�n���9$�`6<��>��E�������xC&~����E�Okb�ɹ>7Ɠqӎ~���`�&i`遼���6��@�^�]$�T��r�҂8��&(s�,��Z�Ao�yq�2<3Lvl���'5ݶ���b<���T�ab׎��nZ���Y�V�>y�3�nJ8�#ޜùwl�xh'�)ɬ��N���D%w���V�N�G7[�j��j�*@�picf�?�iKH%_Opa2���=�89�'���[K���㉉����&ӈd�P�J7z�=	�����C) �C�ko	�(]�Ta3���E<X`��i��]�0�/M����6s�Η��G~G��< �j�5!����U�A#3����50鹁���o�uL왺�)U~�����y�j��H6���h[r�e8������Wf���a��\���k�P!�V=V���� �[7V+�Rt1�f@�0H
!�L���L�<G#C�g���a���i�����VkJ���ǵ��'Sz�|Ϧ��H�q
��K����_����i�s�6Ci�Y�2�1@�ƍid�g�v�`t��&��QOK5cV�A0"�#�'������V����A�R.� ��WM�F�lξp�W.���a�1���$A�£��|#��Y��oȱ��E���/��}H�e���<jJS��*�3��c� �e�x��KG�'�:h���q���K�<M�Λ�B�K{�Qo-YUL!�&�.DU*��Y���L3�HͿT�L֤I����F`4��;s��{�[�v�x	O���'?�k��U�ݠ�@E*I2�)9�P)d����	�v*�C�7M�	�f*^�W�����c�j��c�x�w��~fI�R�)�Ɍ5gᢚ"�a��$�g�@~c�m�j3�|�����,=��	�b�8���}�w&b���D0���7I=`��2 �acf�����~<�'���[�K�G8B����k��V�~/�N� ��
]R�g�,F>�5� ���qrE"�9����VoI���[��!���2	�*�'�袏˹ʧd�@�����Xذ�*�xდ�`]���eL�5]�z�BV�l��c~�����iO�(���ҽQ�f�ֵ����zU�@XBT�����`r]�4���~Ll��%=W��c��g�F���~����&qMOM쮿��|r�H#�;��qe��;�8��9A7T�_o�2���N�̓#�����r�-wC���M�|��b!�Ë��5M��.h��҈��We��c���I(6�c�OX���M�����&��}4�K�f�S�`�
[7B�7@����>r0ՙY��gb�QC��w�ȈS_&�W\s2V��@go�*넖�1��8߁��%�/9���"��'�ٗ�?�@��t�o�'�	��(��Cr.)NO:O'�����5\ww/y�֎�����Nx��	Bb��z� ����]��ʰO�{���|ƺW��T����L� ��(	�܇NR� +A4�N����U�I��~��^6��u&��|�K�x�5������r#v���P��2�ΔM�,Sw�xb���R��ί0�@���k�!��e���e0K���^��~������_�В�"L	��P ycB���w#��GvdP��]NtT�h��М�ll(
�q�+������l"o��֒֔%܂�Fƿ�4/��
ÿ�4��C���2=v�E[=��"�ˊ���� �
`�����Ҵ�}Ө���A<t�>�B5E�u����IԈA*�pp��VOY�����Uf$�,z�rLZ�HJAȃA�c�r^�>6�82+�_H�:x
�M0�ӕV#j��7�p��M]��E��vb¡��l�@�'sKԓ�-!��2��
{�n�U)�Ѥ/q�h���o8@~N4�n������\%A��Vz���}Z�.	��l��<����]񛑍2�k⊕/����$T���F�Kz&���λ3��᤼+CT�*)>uy"ϖ����t��=9	!��ݢ�(�R�����z,5J�L��kO;#�`��8��L����!"���em��5��?'9��N��m��;Veߊ�=)��b/�,{�"�� �<mz��_�d�gO��=���x���2v���v� �C~Z��p��@�3�7���������Q��,?����?CN~�s2�Mԩo���x>��#��nP(����,-d���;��ܭ	7���KDL7��&��#,C�C�X4C\�.����1;@F�VTdmn_�=urt(5�����2�w�
%WI���n�9�ti�h�����#�)��r��h4�!� ��0��y�{�����G��L���6���QG3(��h����J�Iq��݆���:LY"�ۇ�E[�>���9�j��'
� �,�Z�?r�y�ä0��6SDY�ɳN2��k�t���Ca����I��eL<��ݯ����wn�4)Y����M��-r�9{� dSZ�D���r���
ƥ�ĸ��c�_�^䮑�>#M��y��[�k�,���v���a2��ۦįw�&�wvhȂ�/X�'��1t���e�7f�gCi����˃�Y�HLU�!P�����X�� 5���|Ȭq�	e��K��3���f�OjU@��pE\c��*��.��!�B���i���=̌K���60ɤT&3�;�BGt[I��rW9Z�&qE�/{Ѧf�*����]�@�O��y���*F�}���gk�.H>������{&��}�n�0S��L52 ���e*�?I�c~����9�t��x��|����+	��6���.��&mm�)e���^�Rն�n5u����������[Y�"#q3!�c1��bʄ<��� 6	�꾧 O�s�8�ix���[���n���n���bPtl���-T�t�W����GK�H�2\$�0/��?���L\��D�(���v�0�I<Xc�_M��>�WUQgܖT��ѱ`���ـ�	_�e����P�<�����X���p�Ji|��0�.�v�%����Gh<���+�8EL��q��f��zY'����7㧛����}����]��랩�zS�J��i�Ė��