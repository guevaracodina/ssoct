��/  K���D<*J��S���J��S���J��S���J��S���J��S���J��S���J��S���;��o�b?˿�J�eC�J��S������!P7T�Y_"�c�J6�qQ��iQ�����Z:��]ӼPF��+"�N�J6�qQ��J6�qQ��J6�qQ��J6�qQ�^!�t=��+H�Eǋ7=+��	@���;����'��%Ճ�ؿa8�q?*����r�>>7�*m��9Y��d�{Ⱥ��ra�����~f��0(�zފ$0O��1�ljg�w�P�S��Ij�xlP|�gZ.��.�m]	ƞ���{�����薅�#L���*y-w�]����b��Ye���⢵8s%���|߼
�d�g���=[܈uQ��@H��5�+F�-ecȯH5��T��� ���	>^��}V����(_��BD�������abB=]������'ݣ�X�0PW+'�|z��rp$��ρ-��cs1�Ph��Ϸg�~p!ۓ��@�1�_Jz���Uz�(�w1�F���B�șXH#;4ep!!v*!���g�]7~���Onڱ�fǜ��ǽIt��CF)x�es]��M�z ���=��>���i?,�B/R�.��}Բ�p�@�.�S�
)%)���2`萧S����1VCy��@�+O��-��E}m���j�6�S��b;(@��V�(&)~U�Y���k�6�XW�e� T�跤="����{�m:����ie�+:�pW�%�JRz�j>�-H���)X��NcL�5�����b���g#��`ߊ&O0��O�����"�_Zl��H}ꦉ���f%��ڲK�$*�1��N4�X��ť$^N���!Z:c#v��2`萧S������o���1�0�(�3b�4x�����ncst�WC>*��@��f���Ԅ�D�1��.-D)>ƾ~���($�J.���
��'p�@�$���I��m?__� #���P�uorǟD�ui&�%ċ(	q��Ep�/��6�?ʆ�In��tk"3Z"�k�^P��e�G	�S�y�a�\�����Ş4=�-��Ƅ���yM�ꙺi3<�f�D���X���`	SN��r�J��7�8d�������&��J���0�2i#@���%&[?��}	$)wv��I�o��C!T*Y�{'%s��jb�ܳ���7�����������������%������b3�'���Xw�j�7��	��	d��ê����R�wX��W�Px:'0��C�Ό�Z鎬����a�gN�3c!�`�(i3!�`�(i3��6��-G�B$~E��׮�~�b)I��w��,c�A�L'�m��:"�9�2.����T�\ �͌o���F/9
�!�Y`�F����h�7�Gg�����a�O�9� Oag���Ȇ�\�C�l��1J��HI�~|���Fl�	�ȧ��������x	߭��5eqȉ��kz�PՊ(��I�wkGA���G���T�6�ǌ�lAr.��