--megafunction wizard: %Altera SOPC Builder%
--GENERATION: STANDARD
--VERSION: WM1.0


--Legal Notice: (C)2009 Altera Corporation. All rights reserved.  Your
--use of Altera Corporation's design tools, logic functions and other
--software and tools, and its AMPP partner logic functions, and any
--output files any of the foregoing (including device programming or
--simulation files), and any associated documentation or information are
--expressly subject to the terms and conditions of the Altera Program
--License Subscription Agreement or other applicable license agreement,
--including, without limitation, that your use is for the sole purpose
--of programming logic devices manufactured by Altera and sold by Altera
--or its authorized distributors.  Please refer to the applicable
--agreement for further details.


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arbitrator is 
        port (
              -- inputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_read : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reset_n : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_write : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : OUT STD_LOGIC
              );
end entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arbitrator;


architecture europa of NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arbitrator is
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_allgrants :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_allow_new_arb_cycle :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_any_continuerequest :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_counter_enable :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_beginbursttransfer_internal :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_begins_xfer :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_firsttransfer :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_grant_vector :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_in_a_read_cycle :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_in_a_write_cycle :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_master_qreq_vector :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_non_bursting_master_requests :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reg_firsttransfer :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_slavearbiterlockenable :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_unreg_firsttransfer :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waits_for_read :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in :  STD_LOGIC;
                signal shifted_address_to_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer;
    end if;

  end process;

  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in);
  --assign NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa = NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata;
  internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1000000000001000000000000")))) AND pipeline_bridge_m1_chipselect;
  --assign NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa = NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter set values, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_set_values <= std_logic_vector'("001");
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_non_bursting_master_requests mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_any_bursting_master_saved_grant mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_any_bursting_master_saved_grant <= std_logic'('0');
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter_next_value assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_allgrants all slave grants, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_allgrants <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_grant_vector;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer <= NOT ((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waits_for_read OR NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waits_for_write));
  --end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer AND (((NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter arbitration counter enable, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_allgrants)) OR ((end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_non_bursting_master_requests));
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_counter_enable) = '1' then 
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_master_qreq_vector AND end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in)) OR ((end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_non_bursting_master_requests)))) = '1' then 
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_slavearbiterlockenable <= or_reduce(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/in arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_slavearbiterlockenable2 <= or_reduce(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arb_share_counter_next_value);
  --pipeline_bridge/m1 NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/in arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_any_continuerequest at least one master continues requesting, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in <= internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in, which is an e_mux
  pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in <= (internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waits_for_read;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_writedata mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_writedata <= pipeline_bridge_m1_writedata (15 DOWNTO 0);
  --assign NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa = NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket;
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in <= internal_pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in;
  --pipeline_bridge/m1 saved-grant NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/in, which is an e_assign
  pipeline_bridge_m1_saved_grant_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in <= internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in;
  --allow new arb cycle for NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/in, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_master_qreq_vector <= std_logic'('1');
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reset_n assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reset_n <= reset_n;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_firsttransfer first transaction, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_firsttransfer <= A_WE_StdLogic((std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_begins_xfer) = '1'), NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_unreg_firsttransfer, NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reg_firsttransfer);
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_unreg_firsttransfer first transaction, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_unreg_firsttransfer <= NOT ((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_slavearbiterlockenable AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_any_continuerequest));
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_begins_xfer) = '1' then 
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reg_firsttransfer <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_beginbursttransfer_internal <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_begins_xfer;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_read assignment, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_read <= internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_write assignment, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_write <= internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  shifted_address_to_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_address mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_address <= A_EXT (A_SRL(shifted_address_to_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 4);
  --slaveid NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_nativeaddress nativeaddress mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_nativeaddress <= A_EXT (A_SRL(pipeline_bridge_m1_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer;
    end if;

  end process;

  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waits_for_read in a cycle, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waits_for_read <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_in_a_read_cycle AND internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_in_a_read_cycle assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_in_a_read_cycle;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waits_for_write in a cycle, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waits_for_write <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_in_a_write_cycle AND internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_in_a_write_cycle assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_in_a_write_cycle;
  wait_for_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_counter <= std_logic'('0');
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_byteenable byte enable port mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pipeline_bridge_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in <= internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in <= internal_pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in <= internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in;
--synthesis translate_off
    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line, now);
          write(write_line, string'(": "));
          write(write_line, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/in"));
          write(output, write_line.all);
          deallocate (write_line);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_arbitrator is 
        port (
              -- inputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_data_valid_pll_s1 : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1 : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_pll_s1_end_xfer : IN STD_LOGIC;
                 signal pll_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_reset_n : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest : OUT STD_LOGIC
              );
end entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_arbitrator;


architecture europa of NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_arbitrator is
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_last_time :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_run :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write_last_time :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 OR NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_pll_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 OR NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_run <= r_1;
  --optimize select-logic by passing only those address bits which matter.
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/out readdata mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_readdata <= pll_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest <= NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_run;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_reset_n assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave;
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest;
--synthesis translate_off
    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_last_time <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest AND ((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read OR NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write));
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line1 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address /= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_last_time))))) = '1' then 
          write(write_line1, now);
          write(write_line1, string'(": "));
          write(write_line1, string'("NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address did not heed wait!!!"));
          write(output, write_line1.all);
          deallocate (write_line1);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable_last_time <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line2 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable /= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable_last_time))))) = '1' then 
          write(write_line2, now);
          write(write_line2, string'(": "));
          write(write_line2, string'("NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable did not heed wait!!!"));
          write(output, write_line2.all);
          deallocate (write_line2);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_last_time <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line3 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read) /= std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_last_time)))))) = '1' then 
          write(write_line3, now);
          write(write_line3, string'(": "));
          write(write_line3, string'("NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read did not heed wait!!!"));
          write(output, write_line3.all);
          deallocate (write_line3);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write_last_time <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line4 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write) /= std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write_last_time)))))) = '1' then 
          write(write_line4, now);
          write(write_line4, string'(": "));
          write(write_line4, string'("NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write did not heed wait!!!"));
          write(output, write_line4.all);
          deallocate (write_line4);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata_last_time <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line5 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata /= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata_last_time)))) AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write)) = '1' then 
          write(write_line5, now);
          write(write_line5, string'(": "));
          write(write_line5, string'("NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata did not heed wait!!!"));
          write(output, write_line5.all);
          deallocate (write_line5);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arbitrator is 
        port (
              -- inputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_read : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reset_n : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_write : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : OUT STD_LOGIC
              );
end entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arbitrator;


architecture europa of NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arbitrator is
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_allgrants :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_allow_new_arb_cycle :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_any_bursting_master_saved_grant :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_any_continuerequest :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_counter_enable :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_beginbursttransfer_internal :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_begins_xfer :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_firsttransfer :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_grant_vector :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_in_a_read_cycle :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_in_a_write_cycle :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_master_qreq_vector :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_non_bursting_master_requests :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reg_firsttransfer :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_slavearbiterlockenable :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_slavearbiterlockenable2 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_unreg_firsttransfer :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waits_for_read :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in :  STD_LOGIC;
                signal shifted_address_to_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer;
    end if;

  end process;

  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in);
  --assign NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa = NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata;
  internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1000000000001000000100000")))) AND pipeline_bridge_m1_chipselect;
  --assign NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa = NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter set values, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_set_values <= std_logic_vector'("001");
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_non_bursting_master_requests mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_any_bursting_master_saved_grant mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_any_bursting_master_saved_grant <= std_logic'('0');
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter_next_value assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_allgrants all slave grants, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_allgrants <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_grant_vector;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer <= NOT ((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waits_for_read OR NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waits_for_write));
  --end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer AND (((NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter arbitration counter enable, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_counter_enable <= ((end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_allgrants)) OR ((end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_non_bursting_master_requests));
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_counter_enable) = '1' then 
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_master_qreq_vector AND end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in)) OR ((end_xfer_arb_share_counter_term_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_non_bursting_master_requests)))) = '1' then 
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_slavearbiterlockenable <= or_reduce(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/in arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_slavearbiterlockenable2 <= or_reduce(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arb_share_counter_next_value);
  --pipeline_bridge/m1 NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/in arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_any_continuerequest at least one master continues requesting, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in <= internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in, which is an e_mux
  pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in <= (internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waits_for_read;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_writedata mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_writedata <= pipeline_bridge_m1_writedata (15 DOWNTO 0);
  --assign NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa = NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket;
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in <= internal_pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in;
  --pipeline_bridge/m1 saved-grant NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/in, which is an e_assign
  pipeline_bridge_m1_saved_grant_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in <= internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in;
  --allow new arb cycle for NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/in, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_master_qreq_vector <= std_logic'('1');
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reset_n assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reset_n <= reset_n;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_firsttransfer first transaction, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_firsttransfer <= A_WE_StdLogic((std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_begins_xfer) = '1'), NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_unreg_firsttransfer, NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reg_firsttransfer);
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_unreg_firsttransfer first transaction, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_unreg_firsttransfer <= NOT ((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_slavearbiterlockenable AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_any_continuerequest));
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_begins_xfer) = '1' then 
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reg_firsttransfer <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_beginbursttransfer_internal begin burst transfer, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_beginbursttransfer_internal <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_begins_xfer;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_read assignment, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_read <= internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_write assignment, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_write <= internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  shifted_address_to_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_address mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_address <= A_EXT (A_SRL(shifted_address_to_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 4);
  --slaveid NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_nativeaddress nativeaddress mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_nativeaddress <= A_EXT (A_SRL(pipeline_bridge_m1_address_to_slave,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer;
    end if;

  end process;

  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waits_for_read in a cycle, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waits_for_read <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_in_a_read_cycle AND internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_in_a_read_cycle assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_in_a_read_cycle;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waits_for_write in a cycle, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waits_for_write <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_in_a_write_cycle AND internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_in_a_write_cycle assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_in_a_write_cycle;
  wait_for_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_counter <= std_logic'('0');
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_byteenable byte enable port mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pipeline_bridge_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 2);
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in <= internal_pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in <= internal_pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in <= internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in;
--synthesis translate_off
    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/in enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line6 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line6, now);
          write(write_line6, string'(": "));
          write(write_line6, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/in"));
          write(output, write_line6.all);
          deallocate (write_line6);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_arbitrator is 
        port (
              -- inputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_data_valid_tse_pll_s1 : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1 : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal d1_tse_pll_s1_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal tse_pll_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_reset_n : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest : OUT STD_LOGIC
              );
end entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_arbitrator;


architecture europa of NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_arbitrator is
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable_last_time :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_last_time :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_run :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write_last_time :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata_last_time :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001") AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 OR NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_tse_pll_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 OR NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write)))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write)))))))));
  --cascaded wait assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_run <= r_2;
  --optimize select-logic by passing only those address bits which matter.
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/out readdata mux, which is an e_mux
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_readdata <= tse_pll_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest <= NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_run;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_reset_n assignment, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_reset_n <= reset_n;
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave;
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest;
--synthesis translate_off
    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_last_time <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/out waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest AND ((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read OR NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write));
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line7 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address /= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_last_time))))) = '1' then 
          write(write_line7, now);
          write(write_line7, string'(": "));
          write(write_line7, string'("NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address did not heed wait!!!"));
          write(output, write_line7.all);
          deallocate (write_line7);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable_last_time <= std_logic_vector'("00");
      elsif clk'event and clk = '1' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable_last_time <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line8 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable /= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable_last_time))))) = '1' then 
          write(write_line8, now);
          write(write_line8, string'(": "));
          write(write_line8, string'("NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable did not heed wait!!!"));
          write(output, write_line8.all);
          deallocate (write_line8);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_last_time <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line9 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read) /= std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_last_time)))))) = '1' then 
          write(write_line9, now);
          write(write_line9, string'(": "));
          write(write_line9, string'("NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read did not heed wait!!!"));
          write(output, write_line9.all);
          deallocate (write_line9);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write_last_time <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line10 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write) /= std_logic'(NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write_last_time)))))) = '1' then 
          write(write_line10, now);
          write(write_line10, string'(": "));
          write(write_line10, string'("NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write did not heed wait!!!"));
          write(output, write_line10.all);
          deallocate (write_line10);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata_last_time <= std_logic_vector'("0000000000000000");
      elsif clk'event and clk = '1' then
        NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata_last_time <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata;
      end if;

    end process;

    --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line11 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata /= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata_last_time)))) AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write)) = '1' then 
          write(write_line11, now);
          write(write_line11, string'(": "));
          write(write_line11, string'("NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata did not heed wait!!!"));
          write(output, write_line11.all);
          deallocate (write_line11);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity bswap_s1_arbitrator is 
        port (
              -- inputs:
                 signal bswap_s1_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal bswap_s1_select : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal cpu_custom_instruction_master_combo_dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_custom_instruction_master_combo_datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal bswap_s1_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal bswap_s1_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal bswap_s1_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity bswap_s1_arbitrator;


architecture europa of bswap_s1_arbitrator is

begin

  bswap_s1_dataa <= cpu_custom_instruction_master_combo_dataa;
  bswap_s1_datab <= cpu_custom_instruction_master_combo_datab;
  --assign bswap_s1_result_from_sa = bswap_s1_result so that symbol knows where to group signals which may go to master only, which is an e_assign
  bswap_s1_result_from_sa <= bswap_s1_result;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity button_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal button_pio_s1_irq : IN STD_LOGIC;
                 signal button_pio_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal button_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal button_pio_s1_chipselect : OUT STD_LOGIC;
                 signal button_pio_s1_irq_from_sa : OUT STD_LOGIC;
                 signal button_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal button_pio_s1_reset_n : OUT STD_LOGIC;
                 signal button_pio_s1_write_n : OUT STD_LOGIC;
                 signal button_pio_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal d1_button_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_button_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_button_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_button_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_button_pio_s1 : OUT STD_LOGIC
              );
end entity button_pio_s1_arbitrator;


architecture europa of button_pio_s1_arbitrator is
                signal button_pio_s1_allgrants :  STD_LOGIC;
                signal button_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal button_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal button_pio_s1_any_continuerequest :  STD_LOGIC;
                signal button_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal button_pio_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal button_pio_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal button_pio_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal button_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal button_pio_s1_begins_xfer :  STD_LOGIC;
                signal button_pio_s1_end_xfer :  STD_LOGIC;
                signal button_pio_s1_firsttransfer :  STD_LOGIC;
                signal button_pio_s1_grant_vector :  STD_LOGIC;
                signal button_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal button_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal button_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal button_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal button_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal button_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal button_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal button_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal button_pio_s1_waits_for_read :  STD_LOGIC;
                signal button_pio_s1_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_button_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_button_pio_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_button_pio_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_button_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_button_pio_s1 :  STD_LOGIC;
                signal shifted_address_to_button_pio_s1_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_button_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT button_pio_s1_end_xfer;
    end if;

  end process;

  button_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_button_pio_s1);
  --assign button_pio_s1_readdata_from_sa = button_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  button_pio_s1_readdata_from_sa <= button_pio_s1_readdata;
  internal_pipeline_bridge_m1_requests_button_pio_s1 <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000000001000010010000")))) AND pipeline_bridge_m1_chipselect;
  --button_pio_s1_arb_share_counter set values, which is an e_mux
  button_pio_s1_arb_share_set_values <= std_logic_vector'("001");
  --button_pio_s1_non_bursting_master_requests mux, which is an e_mux
  button_pio_s1_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_button_pio_s1;
  --button_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  button_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --button_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  button_pio_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(button_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (button_pio_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(button_pio_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (button_pio_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --button_pio_s1_allgrants all slave grants, which is an e_mux
  button_pio_s1_allgrants <= button_pio_s1_grant_vector;
  --button_pio_s1_end_xfer assignment, which is an e_assign
  button_pio_s1_end_xfer <= NOT ((button_pio_s1_waits_for_read OR button_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_button_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_button_pio_s1 <= button_pio_s1_end_xfer AND (((NOT button_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --button_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  button_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_button_pio_s1 AND button_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_button_pio_s1 AND NOT button_pio_s1_non_bursting_master_requests));
  --button_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      button_pio_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(button_pio_s1_arb_counter_enable) = '1' then 
        button_pio_s1_arb_share_counter <= button_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --button_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      button_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((button_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_button_pio_s1)) OR ((end_xfer_arb_share_counter_term_button_pio_s1 AND NOT button_pio_s1_non_bursting_master_requests)))) = '1' then 
        button_pio_s1_slavearbiterlockenable <= or_reduce(button_pio_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 button_pio/s1 arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= button_pio_s1_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --button_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  button_pio_s1_slavearbiterlockenable2 <= or_reduce(button_pio_s1_arb_share_counter_next_value);
  --pipeline_bridge/m1 button_pio/s1 arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= button_pio_s1_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --button_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  button_pio_s1_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_button_pio_s1 <= internal_pipeline_bridge_m1_requests_button_pio_s1 AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_button_pio_s1, which is an e_mux
  pipeline_bridge_m1_read_data_valid_button_pio_s1 <= (internal_pipeline_bridge_m1_granted_button_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT button_pio_s1_waits_for_read;
  --button_pio_s1_writedata mux, which is an e_mux
  button_pio_s1_writedata <= pipeline_bridge_m1_writedata (3 DOWNTO 0);
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_button_pio_s1 <= internal_pipeline_bridge_m1_qualified_request_button_pio_s1;
  --pipeline_bridge/m1 saved-grant button_pio/s1, which is an e_assign
  pipeline_bridge_m1_saved_grant_button_pio_s1 <= internal_pipeline_bridge_m1_requests_button_pio_s1;
  --allow new arb cycle for button_pio/s1, which is an e_assign
  button_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  button_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  button_pio_s1_master_qreq_vector <= std_logic'('1');
  --button_pio_s1_reset_n assignment, which is an e_assign
  button_pio_s1_reset_n <= reset_n;
  button_pio_s1_chipselect <= internal_pipeline_bridge_m1_granted_button_pio_s1;
  --button_pio_s1_firsttransfer first transaction, which is an e_assign
  button_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(button_pio_s1_begins_xfer) = '1'), button_pio_s1_unreg_firsttransfer, button_pio_s1_reg_firsttransfer);
  --button_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  button_pio_s1_unreg_firsttransfer <= NOT ((button_pio_s1_slavearbiterlockenable AND button_pio_s1_any_continuerequest));
  --button_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      button_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(button_pio_s1_begins_xfer) = '1' then 
        button_pio_s1_reg_firsttransfer <= button_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --button_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  button_pio_s1_beginbursttransfer_internal <= button_pio_s1_begins_xfer;
  --~button_pio_s1_write_n assignment, which is an e_mux
  button_pio_s1_write_n <= NOT ((internal_pipeline_bridge_m1_granted_button_pio_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect))));
  shifted_address_to_button_pio_s1_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --button_pio_s1_address mux, which is an e_mux
  button_pio_s1_address <= A_EXT (A_SRL(shifted_address_to_button_pio_s1_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_button_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_button_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_button_pio_s1_end_xfer <= button_pio_s1_end_xfer;
    end if;

  end process;

  --button_pio_s1_waits_for_read in a cycle, which is an e_mux
  button_pio_s1_waits_for_read <= button_pio_s1_in_a_read_cycle AND button_pio_s1_begins_xfer;
  --button_pio_s1_in_a_read_cycle assignment, which is an e_assign
  button_pio_s1_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_button_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= button_pio_s1_in_a_read_cycle;
  --button_pio_s1_waits_for_write in a cycle, which is an e_mux
  button_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(button_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --button_pio_s1_in_a_write_cycle assignment, which is an e_assign
  button_pio_s1_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_button_pio_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= button_pio_s1_in_a_write_cycle;
  wait_for_button_pio_s1_counter <= std_logic'('0');
  --assign button_pio_s1_irq_from_sa = button_pio_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  button_pio_s1_irq_from_sa <= button_pio_s1_irq;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_button_pio_s1 <= internal_pipeline_bridge_m1_granted_button_pio_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_button_pio_s1 <= internal_pipeline_bridge_m1_qualified_request_button_pio_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_button_pio_s1 <= internal_pipeline_bridge_m1_requests_button_pio_s1;
--synthesis translate_off
    --button_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line12 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_button_pio_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line12, now);
          write(write_line12, string'(": "));
          write(write_line12, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave button_pio/s1"));
          write(output, write_line12.all);
          deallocate (write_line12);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_jtag_debug_module_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_debugaccess : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                 signal cpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_jtag_debug_module_reset : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_write : OUT STD_LOGIC;
                 signal cpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_cpu_jtag_debug_module_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_cpu_jtag_debug_module : OUT STD_LOGIC
              );
end entity cpu_jtag_debug_module_arbitrator;


architecture europa of cpu_jtag_debug_module_arbitrator is
                signal cpu_jtag_debug_module_allgrants :  STD_LOGIC;
                signal cpu_jtag_debug_module_allow_new_arb_cycle :  STD_LOGIC;
                signal cpu_jtag_debug_module_any_bursting_master_saved_grant :  STD_LOGIC;
                signal cpu_jtag_debug_module_any_continuerequest :  STD_LOGIC;
                signal cpu_jtag_debug_module_arb_counter_enable :  STD_LOGIC;
                signal cpu_jtag_debug_module_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal cpu_jtag_debug_module_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal cpu_jtag_debug_module_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal cpu_jtag_debug_module_beginbursttransfer_internal :  STD_LOGIC;
                signal cpu_jtag_debug_module_begins_xfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_firsttransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_grant_vector :  STD_LOGIC;
                signal cpu_jtag_debug_module_in_a_read_cycle :  STD_LOGIC;
                signal cpu_jtag_debug_module_in_a_write_cycle :  STD_LOGIC;
                signal cpu_jtag_debug_module_master_qreq_vector :  STD_LOGIC;
                signal cpu_jtag_debug_module_non_bursting_master_requests :  STD_LOGIC;
                signal cpu_jtag_debug_module_reg_firsttransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_slavearbiterlockenable :  STD_LOGIC;
                signal cpu_jtag_debug_module_slavearbiterlockenable2 :  STD_LOGIC;
                signal cpu_jtag_debug_module_unreg_firsttransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_waits_for_read :  STD_LOGIC;
                signal cpu_jtag_debug_module_waits_for_write :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_cpu_jtag_debug_module :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_cpu_jtag_debug_module :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_cpu_jtag_debug_module :  STD_LOGIC;
                signal shifted_address_to_cpu_jtag_debug_module_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_cpu_jtag_debug_module_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT cpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  cpu_jtag_debug_module_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module);
  --assign cpu_jtag_debug_module_readdata_from_sa = cpu_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_jtag_debug_module_readdata_from_sa <= cpu_jtag_debug_module_readdata;
  internal_pipeline_bridge_m1_requests_cpu_jtag_debug_module <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 11) & std_logic_vector'("00000000000")) = std_logic_vector'("1000000000000000000000000")))) AND pipeline_bridge_m1_chipselect;
  --cpu_jtag_debug_module_arb_share_counter set values, which is an e_mux
  cpu_jtag_debug_module_arb_share_set_values <= std_logic_vector'("001");
  --cpu_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  cpu_jtag_debug_module_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_cpu_jtag_debug_module;
  --cpu_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  cpu_jtag_debug_module_any_bursting_master_saved_grant <= std_logic'('0');
  --cpu_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  cpu_jtag_debug_module_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(cpu_jtag_debug_module_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (cpu_jtag_debug_module_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(cpu_jtag_debug_module_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (cpu_jtag_debug_module_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --cpu_jtag_debug_module_allgrants all slave grants, which is an e_mux
  cpu_jtag_debug_module_allgrants <= cpu_jtag_debug_module_grant_vector;
  --cpu_jtag_debug_module_end_xfer assignment, which is an e_assign
  cpu_jtag_debug_module_end_xfer <= NOT ((cpu_jtag_debug_module_waits_for_read OR cpu_jtag_debug_module_waits_for_write));
  --end_xfer_arb_share_counter_term_cpu_jtag_debug_module arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_cpu_jtag_debug_module <= cpu_jtag_debug_module_end_xfer AND (((NOT cpu_jtag_debug_module_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --cpu_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  cpu_jtag_debug_module_arb_counter_enable <= ((end_xfer_arb_share_counter_term_cpu_jtag_debug_module AND cpu_jtag_debug_module_allgrants)) OR ((end_xfer_arb_share_counter_term_cpu_jtag_debug_module AND NOT cpu_jtag_debug_module_non_bursting_master_requests));
  --cpu_jtag_debug_module_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_jtag_debug_module_arb_counter_enable) = '1' then 
        cpu_jtag_debug_module_arb_share_counter <= cpu_jtag_debug_module_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((cpu_jtag_debug_module_master_qreq_vector AND end_xfer_arb_share_counter_term_cpu_jtag_debug_module)) OR ((end_xfer_arb_share_counter_term_cpu_jtag_debug_module AND NOT cpu_jtag_debug_module_non_bursting_master_requests)))) = '1' then 
        cpu_jtag_debug_module_slavearbiterlockenable <= or_reduce(cpu_jtag_debug_module_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 cpu/jtag_debug_module arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= cpu_jtag_debug_module_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --cpu_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  cpu_jtag_debug_module_slavearbiterlockenable2 <= or_reduce(cpu_jtag_debug_module_arb_share_counter_next_value);
  --pipeline_bridge/m1 cpu/jtag_debug_module arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= cpu_jtag_debug_module_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --cpu_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_assign
  cpu_jtag_debug_module_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module <= internal_pipeline_bridge_m1_requests_cpu_jtag_debug_module AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module, which is an e_mux
  pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module <= (internal_pipeline_bridge_m1_granted_cpu_jtag_debug_module AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT cpu_jtag_debug_module_waits_for_read;
  --cpu_jtag_debug_module_writedata mux, which is an e_mux
  cpu_jtag_debug_module_writedata <= pipeline_bridge_m1_writedata;
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_cpu_jtag_debug_module <= internal_pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;
  --pipeline_bridge/m1 saved-grant cpu/jtag_debug_module, which is an e_assign
  pipeline_bridge_m1_saved_grant_cpu_jtag_debug_module <= internal_pipeline_bridge_m1_requests_cpu_jtag_debug_module;
  --allow new arb cycle for cpu/jtag_debug_module, which is an e_assign
  cpu_jtag_debug_module_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  cpu_jtag_debug_module_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  cpu_jtag_debug_module_master_qreq_vector <= std_logic'('1');
  cpu_jtag_debug_module_begintransfer <= cpu_jtag_debug_module_begins_xfer;
  --~cpu_jtag_debug_module_reset assignment, which is an e_assign
  cpu_jtag_debug_module_reset <= NOT reset_n;
  --assign cpu_jtag_debug_module_resetrequest_from_sa = cpu_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  cpu_jtag_debug_module_resetrequest_from_sa <= cpu_jtag_debug_module_resetrequest;
  cpu_jtag_debug_module_chipselect <= internal_pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  --cpu_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  cpu_jtag_debug_module_firsttransfer <= A_WE_StdLogic((std_logic'(cpu_jtag_debug_module_begins_xfer) = '1'), cpu_jtag_debug_module_unreg_firsttransfer, cpu_jtag_debug_module_reg_firsttransfer);
  --cpu_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  cpu_jtag_debug_module_unreg_firsttransfer <= NOT ((cpu_jtag_debug_module_slavearbiterlockenable AND cpu_jtag_debug_module_any_continuerequest));
  --cpu_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_jtag_debug_module_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(cpu_jtag_debug_module_begins_xfer) = '1' then 
        cpu_jtag_debug_module_reg_firsttransfer <= cpu_jtag_debug_module_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --cpu_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  cpu_jtag_debug_module_beginbursttransfer_internal <= cpu_jtag_debug_module_begins_xfer;
  --cpu_jtag_debug_module_write assignment, which is an e_mux
  cpu_jtag_debug_module_write <= internal_pipeline_bridge_m1_granted_cpu_jtag_debug_module AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  shifted_address_to_cpu_jtag_debug_module_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --cpu_jtag_debug_module_address mux, which is an e_mux
  cpu_jtag_debug_module_address <= A_EXT (A_SRL(shifted_address_to_cpu_jtag_debug_module_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 9);
  --d1_cpu_jtag_debug_module_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_cpu_jtag_debug_module_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_cpu_jtag_debug_module_end_xfer <= cpu_jtag_debug_module_end_xfer;
    end if;

  end process;

  --cpu_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  cpu_jtag_debug_module_waits_for_read <= cpu_jtag_debug_module_in_a_read_cycle AND cpu_jtag_debug_module_begins_xfer;
  --cpu_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  cpu_jtag_debug_module_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_cpu_jtag_debug_module AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= cpu_jtag_debug_module_in_a_read_cycle;
  --cpu_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  cpu_jtag_debug_module_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --cpu_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  cpu_jtag_debug_module_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_cpu_jtag_debug_module AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= cpu_jtag_debug_module_in_a_write_cycle;
  wait_for_cpu_jtag_debug_module_counter <= std_logic'('0');
  --cpu_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  cpu_jtag_debug_module_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_m1_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pipeline_bridge_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --debugaccess mux, which is an e_mux
  cpu_jtag_debug_module_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_m1_granted_cpu_jtag_debug_module)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_cpu_jtag_debug_module <= internal_pipeline_bridge_m1_granted_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module <= internal_pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_cpu_jtag_debug_module <= internal_pipeline_bridge_m1_requests_cpu_jtag_debug_module;
--synthesis translate_off
    --cpu/jtag_debug_module enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line13 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_cpu_jtag_debug_module AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line13, now);
          write(write_line13, string'(": "));
          write(write_line13, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave cpu/jtag_debug_module"));
          write(output, write_line13.all);
          deallocate (write_line13);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity cpu_custom_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal bswap_s1_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal cpu_custom_instruction_master_combo_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal interrupt_vector_interrupt_vector_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal bswap_s1_select : OUT STD_LOGIC;
                 signal cpu_custom_instruction_master_combo_result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_custom_instruction_master_reset_n : OUT STD_LOGIC;
                 signal interrupt_vector_interrupt_vector_select : OUT STD_LOGIC
              );
end entity cpu_custom_instruction_master_arbitrator;


architecture europa of cpu_custom_instruction_master_arbitrator is
                signal internal_bswap_s1_select :  STD_LOGIC;
                signal internal_interrupt_vector_interrupt_vector_select :  STD_LOGIC;

begin

  --cpu_custom_instruction_master_combo_result mux, which is an e_mux
  cpu_custom_instruction_master_combo_result <= ((A_REP(internal_bswap_s1_select, 32) AND bswap_s1_result_from_sa)) OR ((A_REP(internal_interrupt_vector_interrupt_vector_select, 32) AND interrupt_vector_interrupt_vector_result_from_sa));
  --cpu_custom_instruction_master_reset_n local reset_n, which is an e_assign
  cpu_custom_instruction_master_reset_n <= reset_n;
  internal_interrupt_vector_interrupt_vector_select <= to_std_logic((std_logic'(cpu_custom_instruction_master_combo_n(0)) = std_logic'(std_logic'('1'))));
  internal_bswap_s1_select <= to_std_logic((std_logic'(cpu_custom_instruction_master_combo_n(0)) = std_logic'(std_logic'('0'))));
  --vhdl renameroo for output signals
  bswap_s1_select <= internal_bswap_s1_select;
  --vhdl renameroo for output signals
  interrupt_vector_interrupt_vector_select <= internal_interrupt_vector_interrupt_vector_select;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_data_master_arbitrator is 
        port (
              -- inputs:
                 signal button_pio_s1_irq_from_sa : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_granted_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_descriptor_memory_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_ext_ssram_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_packet_memory_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_data_master_granted_tse_mac_control_port : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_ext_ssram_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_packet_memory_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_data_master_qualified_request_tse_mac_control_port : IN STD_LOGIC;
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ext_ssram_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_packet_memory_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_tse_mac_control_port : IN STD_LOGIC;
                 signal cpu_data_master_requests_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_descriptor_memory_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_ext_ssram_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_packet_memory_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_data_master_requests_tse_mac_control_port : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_ddr_sdram_0_s1_end_xfer : IN STD_LOGIC;
                 signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                 signal d1_ext_ssram_bus_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal d1_packet_memory_s1_end_xfer : IN STD_LOGIC;
                 signal d1_pipeline_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal d1_tse_mac_control_port_end_xfer : IN STD_LOGIC;
                 signal ddr_sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ddr_sdram_0_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                 signal descriptor_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal high_res_timer_s1_irq_from_sa : IN STD_LOGIC;
                 signal incoming_ext_ssram_bus_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                 signal packet_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_csr_irq_from_sa : IN STD_LOGIC;
                 signal sgdma_tx_csr_irq_from_sa : IN STD_LOGIC;
                 signal sys_clk_timer_s1_irq_from_sa : IN STD_LOGIC;
                 signal tse_mac_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_control_port_waitrequest_from_sa : IN STD_LOGIC;
                 signal uart1_s1_irq_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_data_master_latency_counter : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_data_master_readdatavalid : OUT STD_LOGIC;
                 signal cpu_data_master_waitrequest : OUT STD_LOGIC
              );
end entity cpu_data_master_arbitrator;


architecture europa of cpu_data_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpu_data_master_address_last_time :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_data_master_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_data_master_is_granted_some_slave :  STD_LOGIC;
                signal cpu_data_master_read_but_no_slave_selected :  STD_LOGIC;
                signal cpu_data_master_read_last_time :  STD_LOGIC;
                signal cpu_data_master_run :  STD_LOGIC;
                signal cpu_data_master_write_last_time :  STD_LOGIC;
                signal cpu_data_master_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_cpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal internal_cpu_data_master_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_cpu_data_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p1_cpu_data_master_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pre_flush_cpu_data_master_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_ddr_sdram_0_s1 OR NOT cpu_data_master_requests_ddr_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_granted_ddr_sdram_0_s1 OR NOT cpu_data_master_qualified_request_ddr_sdram_0_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_ddr_sdram_0_s1 OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ddr_sdram_0_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_ddr_sdram_0_s1 OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ddr_sdram_0_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_descriptor_memory_s1 OR NOT cpu_data_master_requests_descriptor_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_granted_descriptor_memory_s1 OR NOT cpu_data_master_qualified_request_descriptor_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_descriptor_memory_s1 OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_descriptor_memory_s1 OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_data_master_run <= (r_0 AND r_1) AND r_2;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_ext_ssram_s1 OR NOT cpu_data_master_requests_ext_ssram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_granted_ext_ssram_s1 OR NOT cpu_data_master_qualified_request_ext_ssram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_ext_ssram_s1 OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_ext_ssram_s1 OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_packet_memory_s1 OR NOT cpu_data_master_requests_packet_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_packet_memory_s1 OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_packet_memory_s1 OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_pipeline_bridge_s1 OR NOT cpu_data_master_requests_pipeline_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_granted_pipeline_bridge_s1 OR NOT cpu_data_master_qualified_request_pipeline_bridge_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pipeline_bridge_s1 OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pipeline_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_pipeline_bridge_s1 OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pipeline_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_qualified_request_tse_mac_control_port OR NOT cpu_data_master_requests_tse_mac_control_port)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_tse_mac_control_port OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT tse_mac_control_port_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_data_master_qualified_request_tse_mac_control_port OR NOT ((cpu_data_master_read OR cpu_data_master_write)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT tse_mac_control_port_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_data_master_read OR cpu_data_master_write)))))))))));
  --irq assign, which is an e_assign
  cpu_data_master_irq <= Std_Logic_Vector'(A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(button_pio_s1_irq_from_sa) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(high_res_timer_s1_irq_from_sa) & A_ToStdLogicVector(sys_clk_timer_s1_irq_from_sa) & A_ToStdLogicVector(std_logic'('0')) & A_ToStdLogicVector(jtag_uart_avalon_jtag_slave_irq_from_sa) & A_ToStdLogicVector(uart1_s1_irq_from_sa) & A_ToStdLogicVector(sgdma_rx_csr_irq_from_sa) & A_ToStdLogicVector(sgdma_tx_csr_irq_from_sa));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_data_master_address_to_slave <= cpu_data_master_address(27 DOWNTO 0);
  --cpu_data_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_data_master_read_but_no_slave_selected <= (cpu_data_master_read AND cpu_data_master_run) AND NOT cpu_data_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  cpu_data_master_is_granted_some_slave <= ((((cpu_data_master_granted_ddr_sdram_0_s1 OR cpu_data_master_granted_descriptor_memory_s1) OR cpu_data_master_granted_ext_ssram_s1) OR cpu_data_master_granted_packet_memory_s1) OR cpu_data_master_granted_pipeline_bridge_s1) OR cpu_data_master_granted_tse_mac_control_port;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_cpu_data_master_readdatavalid <= (((cpu_data_master_read_data_valid_ddr_sdram_0_s1 OR cpu_data_master_read_data_valid_descriptor_memory_s1) OR cpu_data_master_read_data_valid_ext_ssram_s1) OR cpu_data_master_read_data_valid_packet_memory_s1) OR cpu_data_master_read_data_valid_pipeline_bridge_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  cpu_data_master_readdatavalid <= (((((((((((cpu_data_master_read_but_no_slave_selected OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_but_no_slave_selected) OR pre_flush_cpu_data_master_readdatavalid) OR cpu_data_master_read_data_valid_tse_mac_control_port;
  --cpu/data_master readdata mux, which is an e_mux
  cpu_data_master_readdata <= ((((((A_REP(NOT cpu_data_master_read_data_valid_ddr_sdram_0_s1, 32) OR ddr_sdram_0_s1_readdata_from_sa)) AND ((A_REP(NOT cpu_data_master_read_data_valid_descriptor_memory_s1, 32) OR descriptor_memory_s1_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_read_data_valid_ext_ssram_s1, 32) OR incoming_ext_ssram_bus_data))) AND ((A_REP(NOT cpu_data_master_read_data_valid_packet_memory_s1, 32) OR packet_memory_s1_readdata_from_sa))) AND ((A_REP(NOT cpu_data_master_read_data_valid_pipeline_bridge_s1, 32) OR pipeline_bridge_s1_readdata_from_sa))) AND ((A_REP(NOT ((cpu_data_master_qualified_request_tse_mac_control_port AND cpu_data_master_read)) , 32) OR tse_mac_control_port_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_cpu_data_master_waitrequest <= NOT cpu_data_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_data_master_latency_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      internal_cpu_data_master_latency_counter <= p1_cpu_data_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_cpu_data_master_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((cpu_data_master_run AND cpu_data_master_read))) = '1'), (std_logic_vector'("000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_cpu_data_master_latency_counter)) /= std_logic_vector'("000")), ((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_data_master_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT ((((((std_logic_vector'("00000000000000000000000000000") & (A_REP(cpu_data_master_requests_descriptor_memory_s1, 3))) AND std_logic_vector'("00000000000000000000000000000001"))) OR (((std_logic_vector'("00000000000000000000000000000") & (A_REP(cpu_data_master_requests_ext_ssram_s1, 3))) AND std_logic_vector'("00000000000000000000000000000101")))) OR (((std_logic_vector'("00000000000000000000000000000") & (A_REP(cpu_data_master_requests_packet_memory_s1, 3))) AND std_logic_vector'("00000000000000000000000000000001")))), 3);
  --vhdl renameroo for output signals
  cpu_data_master_address_to_slave <= internal_cpu_data_master_address_to_slave;
  --vhdl renameroo for output signals
  cpu_data_master_latency_counter <= internal_cpu_data_master_latency_counter;
  --vhdl renameroo for output signals
  cpu_data_master_waitrequest <= internal_cpu_data_master_waitrequest;
--synthesis translate_off
    --cpu_data_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_address_last_time <= std_logic_vector'("0000000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_data_master_address_last_time <= cpu_data_master_address;
      end if;

    end process;

    --cpu/data_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpu_data_master_waitrequest AND ((cpu_data_master_read OR cpu_data_master_write));
      end if;

    end process;

    --cpu_data_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line14 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_data_master_address /= cpu_data_master_address_last_time))))) = '1' then 
          write(write_line14, now);
          write(write_line14, string'(": "));
          write(write_line14, string'("cpu_data_master_address did not heed wait!!!"));
          write(output, write_line14.all);
          deallocate (write_line14);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_data_master_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        cpu_data_master_byteenable_last_time <= cpu_data_master_byteenable;
      end if;

    end process;

    --cpu_data_master_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line15 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_data_master_byteenable /= cpu_data_master_byteenable_last_time))))) = '1' then 
          write(write_line15, now);
          write(write_line15, string'(": "));
          write(write_line15, string'("cpu_data_master_byteenable did not heed wait!!!"));
          write(output, write_line15.all);
          deallocate (write_line15);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_data_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_data_master_read_last_time <= cpu_data_master_read;
      end if;

    end process;

    --cpu_data_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line16 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_data_master_read) /= std_logic'(cpu_data_master_read_last_time)))))) = '1' then 
          write(write_line16, now);
          write(write_line16, string'(": "));
          write(write_line16, string'("cpu_data_master_read did not heed wait!!!"));
          write(output, write_line16.all);
          deallocate (write_line16);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_data_master_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_data_master_write_last_time <= cpu_data_master_write;
      end if;

    end process;

    --cpu_data_master_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line17 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_data_master_write) /= std_logic'(cpu_data_master_write_last_time)))))) = '1' then 
          write(write_line17, now);
          write(write_line17, string'(": "));
          write(write_line17, string'("cpu_data_master_write did not heed wait!!!"));
          write(output, write_line17.all);
          deallocate (write_line17);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_data_master_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_data_master_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_data_master_writedata_last_time <= cpu_data_master_writedata;
      end if;

    end process;

    --cpu_data_master_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line18 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((cpu_data_master_writedata /= cpu_data_master_writedata_last_time)))) AND cpu_data_master_write)) = '1' then 
          write(write_line18, now);
          write(write_line18, string'(": "));
          write(write_line18, string'("cpu_data_master_writedata did not heed wait!!!"));
          write(output, write_line18.all);
          deallocate (write_line18);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity cpu_instruction_master_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_instruction_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_instruction_master_granted_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_granted_ext_ssram_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_granted_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_ext_ssram_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_ext_ssram_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_requests_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_requests_ext_ssram_s1 : IN STD_LOGIC;
                 signal cpu_instruction_master_requests_pipeline_bridge_s1 : IN STD_LOGIC;
                 signal d1_ddr_sdram_0_s1_end_xfer : IN STD_LOGIC;
                 signal d1_ext_ssram_bus_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal d1_pipeline_bridge_s1_end_xfer : IN STD_LOGIC;
                 signal ddr_sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ddr_sdram_0_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                 signal incoming_ext_ssram_bus_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                 signal cpu_instruction_master_waitrequest : OUT STD_LOGIC
              );
end entity cpu_instruction_master_arbitrator;


architecture europa of cpu_instruction_master_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal cpu_instruction_master_address_last_time :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_instruction_master_is_granted_some_slave :  STD_LOGIC;
                signal cpu_instruction_master_read_but_no_slave_selected :  STD_LOGIC;
                signal cpu_instruction_master_read_last_time :  STD_LOGIC;
                signal cpu_instruction_master_run :  STD_LOGIC;
                signal internal_cpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal internal_cpu_instruction_master_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_cpu_instruction_master_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p1_cpu_instruction_master_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pre_flush_cpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_qualified_request_ddr_sdram_0_s1 OR NOT cpu_instruction_master_requests_ddr_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_granted_ddr_sdram_0_s1 OR NOT cpu_instruction_master_qualified_request_ddr_sdram_0_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_instruction_master_qualified_request_ddr_sdram_0_s1 OR NOT (cpu_instruction_master_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ddr_sdram_0_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_read))))))))));
  --cascaded wait assignment, which is an e_assign
  cpu_instruction_master_run <= r_0 AND r_1;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_qualified_request_ext_ssram_s1 OR NOT cpu_instruction_master_requests_ext_ssram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_granted_ext_ssram_s1 OR NOT cpu_instruction_master_qualified_request_ext_ssram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_instruction_master_qualified_request_ext_ssram_s1 OR NOT (cpu_instruction_master_read))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_read))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_qualified_request_pipeline_bridge_s1 OR NOT cpu_instruction_master_requests_pipeline_bridge_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((cpu_instruction_master_granted_pipeline_bridge_s1 OR NOT cpu_instruction_master_qualified_request_pipeline_bridge_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT cpu_instruction_master_qualified_request_pipeline_bridge_s1 OR NOT (cpu_instruction_master_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT pipeline_bridge_s1_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((cpu_instruction_master_read))))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_cpu_instruction_master_address_to_slave <= cpu_instruction_master_address(27 DOWNTO 0);
  --cpu_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_instruction_master_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_instruction_master_read_but_no_slave_selected <= (cpu_instruction_master_read AND cpu_instruction_master_run) AND NOT cpu_instruction_master_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  cpu_instruction_master_is_granted_some_slave <= (cpu_instruction_master_granted_ddr_sdram_0_s1 OR cpu_instruction_master_granted_ext_ssram_s1) OR cpu_instruction_master_granted_pipeline_bridge_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_cpu_instruction_master_readdatavalid <= (cpu_instruction_master_read_data_valid_ddr_sdram_0_s1 OR cpu_instruction_master_read_data_valid_ext_ssram_s1) OR cpu_instruction_master_read_data_valid_pipeline_bridge_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  cpu_instruction_master_readdatavalid <= ((((cpu_instruction_master_read_but_no_slave_selected OR pre_flush_cpu_instruction_master_readdatavalid) OR cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_cpu_instruction_master_readdatavalid) OR cpu_instruction_master_read_but_no_slave_selected) OR pre_flush_cpu_instruction_master_readdatavalid;
  --cpu/instruction_master readdata mux, which is an e_mux
  cpu_instruction_master_readdata <= (((A_REP(NOT cpu_instruction_master_read_data_valid_ddr_sdram_0_s1, 32) OR ddr_sdram_0_s1_readdata_from_sa)) AND ((A_REP(NOT cpu_instruction_master_read_data_valid_ext_ssram_s1, 32) OR incoming_ext_ssram_bus_data))) AND ((A_REP(NOT cpu_instruction_master_read_data_valid_pipeline_bridge_s1, 32) OR pipeline_bridge_s1_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_cpu_instruction_master_waitrequest <= NOT cpu_instruction_master_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_cpu_instruction_master_latency_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      internal_cpu_instruction_master_latency_counter <= p1_cpu_instruction_master_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_cpu_instruction_master_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((cpu_instruction_master_run AND cpu_instruction_master_read))) = '1'), (std_logic_vector'("000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_cpu_instruction_master_latency_counter)) /= std_logic_vector'("000")), ((std_logic_vector'("000000000000000000000000000000") & (internal_cpu_instruction_master_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (A_REP(cpu_instruction_master_requests_ext_ssram_s1, 3))) AND std_logic_vector'("00000000000000000000000000000101")), 3);
  --vhdl renameroo for output signals
  cpu_instruction_master_address_to_slave <= internal_cpu_instruction_master_address_to_slave;
  --vhdl renameroo for output signals
  cpu_instruction_master_latency_counter <= internal_cpu_instruction_master_latency_counter;
  --vhdl renameroo for output signals
  cpu_instruction_master_waitrequest <= internal_cpu_instruction_master_waitrequest;
--synthesis translate_off
    --cpu_instruction_master_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_instruction_master_address_last_time <= std_logic_vector'("0000000000000000000000000000");
      elsif clk'event and clk = '1' then
        cpu_instruction_master_address_last_time <= cpu_instruction_master_address;
      end if;

    end process;

    --cpu/instruction_master waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_cpu_instruction_master_waitrequest AND (cpu_instruction_master_read);
      end if;

    end process;

    --cpu_instruction_master_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line19 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((cpu_instruction_master_address /= cpu_instruction_master_address_last_time))))) = '1' then 
          write(write_line19, now);
          write(write_line19, string'(": "));
          write(write_line19, string'("cpu_instruction_master_address did not heed wait!!!"));
          write(output, write_line19.all);
          deallocate (write_line19);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --cpu_instruction_master_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        cpu_instruction_master_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        cpu_instruction_master_read_last_time <= cpu_instruction_master_read;
      end if;

    end process;

    --cpu_instruction_master_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line20 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(cpu_instruction_master_read) /= std_logic'(cpu_instruction_master_read_last_time)))))) = '1' then 
          write(write_line20, now);
          write(write_line20, string'(": "));
          write(write_line20, string'("cpu_instruction_master_read did not heed wait!!!"));
          write(output, write_line20.all);
          deallocate (write_line20);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_ddr_sdram_0_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_ddr_sdram_0_s1_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_ddr_sdram_0_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_15;
  empty <= NOT(full_0);
  full_16 <= std_logic'('0');
  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 6);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 6);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 6);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_instruction_master_to_ddr_sdram_0_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_instruction_master_to_ddr_sdram_0_s1_module;


architecture europa of rdv_fifo_for_cpu_instruction_master_to_ddr_sdram_0_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_15;
  empty <= NOT(full_0);
  full_16 <= std_logic'('0');
  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 6);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 6);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 6);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_sgdma_tx_m_read_to_ddr_sdram_0_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_sgdma_tx_m_read_to_ddr_sdram_0_s1_module;


architecture europa of rdv_fifo_for_sgdma_tx_m_read_to_ddr_sdram_0_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_10 :  STD_LOGIC;
                signal full_11 :  STD_LOGIC;
                signal full_12 :  STD_LOGIC;
                signal full_13 :  STD_LOGIC;
                signal full_14 :  STD_LOGIC;
                signal full_15 :  STD_LOGIC;
                signal full_16 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal full_6 :  STD_LOGIC;
                signal full_7 :  STD_LOGIC;
                signal full_8 :  STD_LOGIC;
                signal full_9 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p10_full_10 :  STD_LOGIC;
                signal p10_stage_10 :  STD_LOGIC;
                signal p11_full_11 :  STD_LOGIC;
                signal p11_stage_11 :  STD_LOGIC;
                signal p12_full_12 :  STD_LOGIC;
                signal p12_stage_12 :  STD_LOGIC;
                signal p13_full_13 :  STD_LOGIC;
                signal p13_stage_13 :  STD_LOGIC;
                signal p14_full_14 :  STD_LOGIC;
                signal p14_stage_14 :  STD_LOGIC;
                signal p15_full_15 :  STD_LOGIC;
                signal p15_stage_15 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal p5_full_5 :  STD_LOGIC;
                signal p5_stage_5 :  STD_LOGIC;
                signal p6_full_6 :  STD_LOGIC;
                signal p6_stage_6 :  STD_LOGIC;
                signal p7_full_7 :  STD_LOGIC;
                signal p7_stage_7 :  STD_LOGIC;
                signal p8_full_8 :  STD_LOGIC;
                signal p8_stage_8 :  STD_LOGIC;
                signal p9_full_9 :  STD_LOGIC;
                signal p9_stage_9 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_10 :  STD_LOGIC;
                signal stage_11 :  STD_LOGIC;
                signal stage_12 :  STD_LOGIC;
                signal stage_13 :  STD_LOGIC;
                signal stage_14 :  STD_LOGIC;
                signal stage_15 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal stage_5 :  STD_LOGIC;
                signal stage_6 :  STD_LOGIC;
                signal stage_7 :  STD_LOGIC;
                signal stage_8 :  STD_LOGIC;
                signal stage_9 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (5 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_15;
  empty <= NOT(full_0);
  full_16 <= std_logic'('0');
  --data_15, which is an e_mux
  p15_stage_15 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_16 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_15))))) = '1' then 
        if std_logic'(((sync_reset AND full_15) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_16))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_15 <= std_logic'('0');
        else
          stage_15 <= p15_stage_15;
        end if;
      end if;
    end if;

  end process;

  --control_15, which is an e_mux
  p15_full_15 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_15, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_15 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_15 <= std_logic'('0');
        else
          full_15 <= p15_full_15;
        end if;
      end if;
    end if;

  end process;

  --data_14, which is an e_mux
  p14_stage_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_15 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_15);
  --data_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_14))))) = '1' then 
        if std_logic'(((sync_reset AND full_14) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_15))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_14 <= std_logic'('0');
        else
          stage_14 <= p14_stage_14;
        end if;
      end if;
    end if;

  end process;

  --control_14, which is an e_mux
  p14_full_14 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_13, full_15);
  --control_reg_14, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_14 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_14 <= std_logic'('0');
        else
          full_14 <= p14_full_14;
        end if;
      end if;
    end if;

  end process;

  --data_13, which is an e_mux
  p13_stage_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_14 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_14);
  --data_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_13))))) = '1' then 
        if std_logic'(((sync_reset AND full_13) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_14))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_13 <= std_logic'('0');
        else
          stage_13 <= p13_stage_13;
        end if;
      end if;
    end if;

  end process;

  --control_13, which is an e_mux
  p13_full_13 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_12, full_14);
  --control_reg_13, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_13 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_13 <= std_logic'('0');
        else
          full_13 <= p13_full_13;
        end if;
      end if;
    end if;

  end process;

  --data_12, which is an e_mux
  p12_stage_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_13 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_13);
  --data_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_12))))) = '1' then 
        if std_logic'(((sync_reset AND full_12) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_13))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_12 <= std_logic'('0');
        else
          stage_12 <= p12_stage_12;
        end if;
      end if;
    end if;

  end process;

  --control_12, which is an e_mux
  p12_full_12 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_11, full_13);
  --control_reg_12, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_12 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_12 <= std_logic'('0');
        else
          full_12 <= p12_full_12;
        end if;
      end if;
    end if;

  end process;

  --data_11, which is an e_mux
  p11_stage_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_12 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_12);
  --data_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_11))))) = '1' then 
        if std_logic'(((sync_reset AND full_11) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_12))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_11 <= std_logic'('0');
        else
          stage_11 <= p11_stage_11;
        end if;
      end if;
    end if;

  end process;

  --control_11, which is an e_mux
  p11_full_11 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_10, full_12);
  --control_reg_11, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_11 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_11 <= std_logic'('0');
        else
          full_11 <= p11_full_11;
        end if;
      end if;
    end if;

  end process;

  --data_10, which is an e_mux
  p10_stage_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_11 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_11);
  --data_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_10))))) = '1' then 
        if std_logic'(((sync_reset AND full_10) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_11))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_10 <= std_logic'('0');
        else
          stage_10 <= p10_stage_10;
        end if;
      end if;
    end if;

  end process;

  --control_10, which is an e_mux
  p10_full_10 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_9, full_11);
  --control_reg_10, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_10 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_10 <= std_logic'('0');
        else
          full_10 <= p10_full_10;
        end if;
      end if;
    end if;

  end process;

  --data_9, which is an e_mux
  p9_stage_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_10 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_10);
  --data_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_9))))) = '1' then 
        if std_logic'(((sync_reset AND full_9) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_10))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_9 <= std_logic'('0');
        else
          stage_9 <= p9_stage_9;
        end if;
      end if;
    end if;

  end process;

  --control_9, which is an e_mux
  p9_full_9 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_8, full_10);
  --control_reg_9, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_9 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_9 <= std_logic'('0');
        else
          full_9 <= p9_full_9;
        end if;
      end if;
    end if;

  end process;

  --data_8, which is an e_mux
  p8_stage_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_9 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_9);
  --data_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_8))))) = '1' then 
        if std_logic'(((sync_reset AND full_8) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_9))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_8 <= std_logic'('0');
        else
          stage_8 <= p8_stage_8;
        end if;
      end if;
    end if;

  end process;

  --control_8, which is an e_mux
  p8_full_8 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_7, full_9);
  --control_reg_8, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_8 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_8 <= std_logic'('0');
        else
          full_8 <= p8_full_8;
        end if;
      end if;
    end if;

  end process;

  --data_7, which is an e_mux
  p7_stage_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_8 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_8);
  --data_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_7))))) = '1' then 
        if std_logic'(((sync_reset AND full_7) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_8))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_7 <= std_logic'('0');
        else
          stage_7 <= p7_stage_7;
        end if;
      end if;
    end if;

  end process;

  --control_7, which is an e_mux
  p7_full_7 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_6, full_8);
  --control_reg_7, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_7 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_7 <= std_logic'('0');
        else
          full_7 <= p7_full_7;
        end if;
      end if;
    end if;

  end process;

  --data_6, which is an e_mux
  p6_stage_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_7 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_7);
  --data_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_6))))) = '1' then 
        if std_logic'(((sync_reset AND full_6) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_7))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_6 <= std_logic'('0');
        else
          stage_6 <= p6_stage_6;
        end if;
      end if;
    end if;

  end process;

  --control_6, which is an e_mux
  p6_full_6 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_5, full_7);
  --control_reg_6, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_6 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_6 <= std_logic'('0');
        else
          full_6 <= p6_full_6;
        end if;
      end if;
    end if;

  end process;

  --data_5, which is an e_mux
  p5_stage_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_6 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_6);
  --data_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_5))))) = '1' then 
        if std_logic'(((sync_reset AND full_5) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_6))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_5 <= std_logic'('0');
        else
          stage_5 <= p5_stage_5;
        end if;
      end if;
    end if;

  end process;

  --control_5, which is an e_mux
  p5_full_5 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_4, full_6);
  --control_reg_5, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_5 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_5 <= std_logic'('0');
        else
          full_5 <= p5_full_5;
        end if;
      end if;
    end if;

  end process;

  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_5);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_3, full_5);
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 6);
  one_count_minus_one <= A_EXT (((std_logic_vector'("000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 6);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("00000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("00000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 6);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ddr_sdram_0_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal ddr_sdram_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ddr_sdram_0_s1_readdatavalid : IN STD_LOGIC;
                 signal ddr_sdram_0_s1_waitrequest_n : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_m_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal sgdma_rx_m_write_write : IN STD_LOGIC;
                 signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal sgdma_tx_m_read_read : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_granted_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_instruction_master_requests_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal d1_ddr_sdram_0_s1_end_xfer : OUT STD_LOGIC;
                 signal ddr_sdram_0_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal ddr_sdram_0_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal ddr_sdram_0_s1_read : OUT STD_LOGIC;
                 signal ddr_sdram_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ddr_sdram_0_s1_reset_n : OUT STD_LOGIC;
                 signal ddr_sdram_0_s1_waitrequest_n_from_sa : OUT STD_LOGIC;
                 signal ddr_sdram_0_s1_write : OUT STD_LOGIC;
                 signal ddr_sdram_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_m_write_granted_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_m_write_requests_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_granted_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_requests_ddr_sdram_0_s1 : OUT STD_LOGIC
              );
end entity ddr_sdram_0_s1_arbitrator;


architecture europa of ddr_sdram_0_s1_arbitrator is
component rdv_fifo_for_cpu_data_master_to_ddr_sdram_0_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_ddr_sdram_0_s1_module;

component rdv_fifo_for_cpu_instruction_master_to_ddr_sdram_0_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_instruction_master_to_ddr_sdram_0_s1_module;

component rdv_fifo_for_sgdma_tx_m_read_to_ddr_sdram_0_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_sgdma_tx_m_read_to_ddr_sdram_0_s1_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_data_master_saved_grant_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_empty_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_output_from_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_instruction_master_saved_grant_ddr_sdram_0_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal ddr_sdram_0_s1_allgrants :  STD_LOGIC;
                signal ddr_sdram_0_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal ddr_sdram_0_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal ddr_sdram_0_s1_any_continuerequest :  STD_LOGIC;
                signal ddr_sdram_0_s1_arb_addend :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_0_s1_arb_counter_enable :  STD_LOGIC;
                signal ddr_sdram_0_s1_arb_share_counter :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_0_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_0_s1_arb_share_set_values :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_0_s1_arb_winner :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_0_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal ddr_sdram_0_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal ddr_sdram_0_s1_begins_xfer :  STD_LOGIC;
                signal ddr_sdram_0_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal ddr_sdram_0_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_0_s1_end_xfer :  STD_LOGIC;
                signal ddr_sdram_0_s1_firsttransfer :  STD_LOGIC;
                signal ddr_sdram_0_s1_grant_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_0_s1_in_a_read_cycle :  STD_LOGIC;
                signal ddr_sdram_0_s1_in_a_write_cycle :  STD_LOGIC;
                signal ddr_sdram_0_s1_master_qreq_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_0_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal ddr_sdram_0_s1_non_bursting_master_requests :  STD_LOGIC;
                signal ddr_sdram_0_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal ddr_sdram_0_s1_reg_firsttransfer :  STD_LOGIC;
                signal ddr_sdram_0_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_0_s1_slavearbiterlockenable :  STD_LOGIC;
                signal ddr_sdram_0_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal ddr_sdram_0_s1_unreg_firsttransfer :  STD_LOGIC;
                signal ddr_sdram_0_s1_waits_for_read :  STD_LOGIC;
                signal ddr_sdram_0_s1_waits_for_write :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_ddr_sdram_0_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_cpu_instruction_master_granted_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_cpu_instruction_master_qualified_request_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_cpu_instruction_master_requests_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_ddr_sdram_0_s1_waitrequest_n_from_sa :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_granted_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_granted_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1 :  STD_LOGIC;
                signal last_cycle_cpu_data_master_granted_slave_ddr_sdram_0_s1 :  STD_LOGIC;
                signal last_cycle_cpu_instruction_master_granted_slave_ddr_sdram_0_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_rx_m_write_granted_slave_ddr_sdram_0_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_tx_m_read_granted_slave_ddr_sdram_0_s1 :  STD_LOGIC;
                signal module_input :  STD_LOGIC;
                signal module_input1 :  STD_LOGIC;
                signal module_input2 :  STD_LOGIC;
                signal module_input3 :  STD_LOGIC;
                signal module_input4 :  STD_LOGIC;
                signal module_input5 :  STD_LOGIC;
                signal module_input6 :  STD_LOGIC;
                signal module_input7 :  STD_LOGIC;
                signal module_input8 :  STD_LOGIC;
                signal sgdma_rx_m_write_arbiterlock :  STD_LOGIC;
                signal sgdma_rx_m_write_arbiterlock2 :  STD_LOGIC;
                signal sgdma_rx_m_write_continuerequest :  STD_LOGIC;
                signal sgdma_rx_m_write_saved_grant_ddr_sdram_0_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_arbiterlock :  STD_LOGIC;
                signal sgdma_tx_m_read_arbiterlock2 :  STD_LOGIC;
                signal sgdma_tx_m_read_continuerequest :  STD_LOGIC;
                signal sgdma_tx_m_read_rdv_fifo_empty_ddr_sdram_0_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_rdv_fifo_output_from_ddr_sdram_0_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_saved_grant_ddr_sdram_0_s1 :  STD_LOGIC;
                signal shifted_address_to_ddr_sdram_0_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal shifted_address_to_ddr_sdram_0_s1_from_cpu_instruction_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal shifted_address_to_ddr_sdram_0_s1_from_sgdma_rx_m_write :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_ddr_sdram_0_s1_from_sgdma_tx_m_read :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal wait_for_ddr_sdram_0_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT ddr_sdram_0_s1_end_xfer;
    end if;

  end process;

  ddr_sdram_0_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((((internal_cpu_data_master_qualified_request_ddr_sdram_0_s1 OR internal_cpu_instruction_master_qualified_request_ddr_sdram_0_s1) OR internal_sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1) OR internal_sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1));
  --assign ddr_sdram_0_s1_readdata_from_sa = ddr_sdram_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  ddr_sdram_0_s1_readdata_from_sa <= ddr_sdram_0_s1_readdata;
  internal_cpu_data_master_requests_ddr_sdram_0_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(27 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("0010000000000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign ddr_sdram_0_s1_waitrequest_n_from_sa = ddr_sdram_0_s1_waitrequest_n so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_ddr_sdram_0_s1_waitrequest_n_from_sa <= ddr_sdram_0_s1_waitrequest_n;
  --assign ddr_sdram_0_s1_readdatavalid_from_sa = ddr_sdram_0_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  ddr_sdram_0_s1_readdatavalid_from_sa <= ddr_sdram_0_s1_readdatavalid;
  --ddr_sdram_0_s1_arb_share_counter set values, which is an e_mux
  ddr_sdram_0_s1_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ddr_sdram_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_ddr_sdram_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ddr_sdram_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_ddr_sdram_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ddr_sdram_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_ddr_sdram_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ddr_sdram_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_ddr_sdram_0_s1)) = '1'), std_logic_vector'("00000000000000000000000000001000"), std_logic_vector'("00000000000000000000000000000001"))))))))), 4);
  --ddr_sdram_0_s1_non_bursting_master_requests mux, which is an e_mux
  ddr_sdram_0_s1_non_bursting_master_requests <= ((((((((((((((internal_cpu_data_master_requests_ddr_sdram_0_s1 OR internal_cpu_instruction_master_requests_ddr_sdram_0_s1) OR internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1) OR internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1) OR internal_cpu_data_master_requests_ddr_sdram_0_s1) OR internal_cpu_instruction_master_requests_ddr_sdram_0_s1) OR internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1) OR internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1) OR internal_cpu_data_master_requests_ddr_sdram_0_s1) OR internal_cpu_instruction_master_requests_ddr_sdram_0_s1) OR internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1) OR internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1) OR internal_cpu_data_master_requests_ddr_sdram_0_s1) OR internal_cpu_instruction_master_requests_ddr_sdram_0_s1) OR internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1) OR internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1;
  --ddr_sdram_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  ddr_sdram_0_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --ddr_sdram_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  ddr_sdram_0_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(ddr_sdram_0_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (ddr_sdram_0_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(ddr_sdram_0_s1_arb_share_counter)) = '1'), (((std_logic_vector'("00000000000000000000000000000") & (ddr_sdram_0_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 4);
  --ddr_sdram_0_s1_allgrants all slave grants, which is an e_mux
  ddr_sdram_0_s1_allgrants <= (((((((((((((((or_reduce(ddr_sdram_0_s1_grant_vector)) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector))) OR (or_reduce(ddr_sdram_0_s1_grant_vector));
  --ddr_sdram_0_s1_end_xfer assignment, which is an e_assign
  ddr_sdram_0_s1_end_xfer <= NOT ((ddr_sdram_0_s1_waits_for_read OR ddr_sdram_0_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_ddr_sdram_0_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_ddr_sdram_0_s1 <= ddr_sdram_0_s1_end_xfer AND (((NOT ddr_sdram_0_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --ddr_sdram_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  ddr_sdram_0_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_ddr_sdram_0_s1 AND ddr_sdram_0_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_ddr_sdram_0_s1 AND NOT ddr_sdram_0_s1_non_bursting_master_requests));
  --ddr_sdram_0_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ddr_sdram_0_s1_arb_share_counter <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(ddr_sdram_0_s1_arb_counter_enable) = '1' then 
        ddr_sdram_0_s1_arb_share_counter <= ddr_sdram_0_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ddr_sdram_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ddr_sdram_0_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(ddr_sdram_0_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_ddr_sdram_0_s1)) OR ((end_xfer_arb_share_counter_term_ddr_sdram_0_s1 AND NOT ddr_sdram_0_s1_non_bursting_master_requests)))) = '1' then 
        ddr_sdram_0_s1_slavearbiterlockenable <= or_reduce(ddr_sdram_0_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --cpu/data_master ddr_sdram_0/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= ddr_sdram_0_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --ddr_sdram_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  ddr_sdram_0_s1_slavearbiterlockenable2 <= or_reduce(ddr_sdram_0_s1_arb_share_counter_next_value);
  --cpu/data_master ddr_sdram_0/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= ddr_sdram_0_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --cpu/instruction_master ddr_sdram_0/s1 arbiterlock, which is an e_assign
  cpu_instruction_master_arbiterlock <= ddr_sdram_0_s1_slavearbiterlockenable AND cpu_instruction_master_continuerequest;
  --cpu/instruction_master ddr_sdram_0/s1 arbiterlock2, which is an e_assign
  cpu_instruction_master_arbiterlock2 <= ddr_sdram_0_s1_slavearbiterlockenable2 AND cpu_instruction_master_continuerequest;
  --cpu/instruction_master granted ddr_sdram_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_instruction_master_granted_slave_ddr_sdram_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_instruction_master_granted_slave_ddr_sdram_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_instruction_master_saved_grant_ddr_sdram_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((ddr_sdram_0_s1_arbitration_holdoff_internal OR NOT internal_cpu_instruction_master_requests_ddr_sdram_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_instruction_master_granted_slave_ddr_sdram_0_s1))))));
    end if;

  end process;

  --cpu_instruction_master_continuerequest continued request, which is an e_mux
  cpu_instruction_master_continuerequest <= (((last_cycle_cpu_instruction_master_granted_slave_ddr_sdram_0_s1 AND internal_cpu_instruction_master_requests_ddr_sdram_0_s1)) OR ((last_cycle_cpu_instruction_master_granted_slave_ddr_sdram_0_s1 AND internal_cpu_instruction_master_requests_ddr_sdram_0_s1))) OR ((last_cycle_cpu_instruction_master_granted_slave_ddr_sdram_0_s1 AND internal_cpu_instruction_master_requests_ddr_sdram_0_s1));
  --ddr_sdram_0_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  ddr_sdram_0_s1_any_continuerequest <= ((((((((((cpu_instruction_master_continuerequest OR sgdma_rx_m_write_continuerequest) OR sgdma_tx_m_read_continuerequest) OR cpu_data_master_continuerequest) OR sgdma_rx_m_write_continuerequest) OR sgdma_tx_m_read_continuerequest) OR cpu_data_master_continuerequest) OR cpu_instruction_master_continuerequest) OR sgdma_tx_m_read_continuerequest) OR cpu_data_master_continuerequest) OR cpu_instruction_master_continuerequest) OR sgdma_rx_m_write_continuerequest;
  --sgdma_rx/m_write ddr_sdram_0/s1 arbiterlock, which is an e_assign
  sgdma_rx_m_write_arbiterlock <= ddr_sdram_0_s1_slavearbiterlockenable AND sgdma_rx_m_write_continuerequest;
  --sgdma_rx/m_write ddr_sdram_0/s1 arbiterlock2, which is an e_assign
  sgdma_rx_m_write_arbiterlock2 <= ddr_sdram_0_s1_slavearbiterlockenable2 AND sgdma_rx_m_write_continuerequest;
  --sgdma_rx/m_write granted ddr_sdram_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_rx_m_write_granted_slave_ddr_sdram_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_rx_m_write_granted_slave_ddr_sdram_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_rx_m_write_saved_grant_ddr_sdram_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((ddr_sdram_0_s1_arbitration_holdoff_internal OR NOT internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_rx_m_write_granted_slave_ddr_sdram_0_s1))))));
    end if;

  end process;

  --sgdma_rx_m_write_continuerequest continued request, which is an e_mux
  sgdma_rx_m_write_continuerequest <= (((last_cycle_sgdma_rx_m_write_granted_slave_ddr_sdram_0_s1 AND internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1)) OR ((last_cycle_sgdma_rx_m_write_granted_slave_ddr_sdram_0_s1 AND internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1))) OR ((last_cycle_sgdma_rx_m_write_granted_slave_ddr_sdram_0_s1 AND internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1));
  --sgdma_tx/m_read ddr_sdram_0/s1 arbiterlock, which is an e_assign
  sgdma_tx_m_read_arbiterlock <= ddr_sdram_0_s1_slavearbiterlockenable AND sgdma_tx_m_read_continuerequest;
  --sgdma_tx/m_read ddr_sdram_0/s1 arbiterlock2, which is an e_assign
  sgdma_tx_m_read_arbiterlock2 <= ddr_sdram_0_s1_slavearbiterlockenable2 AND sgdma_tx_m_read_continuerequest;
  --sgdma_tx/m_read granted ddr_sdram_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_tx_m_read_granted_slave_ddr_sdram_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_tx_m_read_granted_slave_ddr_sdram_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_tx_m_read_saved_grant_ddr_sdram_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((ddr_sdram_0_s1_arbitration_holdoff_internal OR NOT internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_tx_m_read_granted_slave_ddr_sdram_0_s1))))));
    end if;

  end process;

  --sgdma_tx_m_read_continuerequest continued request, which is an e_mux
  sgdma_tx_m_read_continuerequest <= (((last_cycle_sgdma_tx_m_read_granted_slave_ddr_sdram_0_s1 AND internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1)) OR ((last_cycle_sgdma_tx_m_read_granted_slave_ddr_sdram_0_s1 AND internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1))) OR ((last_cycle_sgdma_tx_m_read_granted_slave_ddr_sdram_0_s1 AND internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1));
  internal_cpu_data_master_qualified_request_ddr_sdram_0_s1 <= internal_cpu_data_master_requests_ddr_sdram_0_s1 AND NOT ((((((cpu_data_master_read AND ((to_std_logic(((((std_logic_vector'("00000000000000000000000000000") & (cpu_data_master_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("00000000000000000000000000000") & (cpu_data_master_latency_counter)))))) OR (cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register))))) OR cpu_instruction_master_arbiterlock) OR sgdma_rx_m_write_arbiterlock) OR sgdma_tx_m_read_arbiterlock));
  --unique name for ddr_sdram_0_s1_move_on_to_next_transaction, which is an e_assign
  ddr_sdram_0_s1_move_on_to_next_transaction <= ddr_sdram_0_s1_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_ddr_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_ddr_sdram_0_s1 : rdv_fifo_for_cpu_data_master_to_ddr_sdram_0_s1_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_ddr_sdram_0_s1,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_ddr_sdram_0_s1,
      full => open,
      clear_fifo => module_input,
      clk => clk,
      data_in => internal_cpu_data_master_granted_ddr_sdram_0_s1,
      read => ddr_sdram_0_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input1,
      write => module_input2
    );

  module_input <= std_logic'('0');
  module_input1 <= std_logic'('0');
  module_input2 <= in_a_read_cycle AND NOT ddr_sdram_0_s1_waits_for_read;

  cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register <= NOT cpu_data_master_rdv_fifo_empty_ddr_sdram_0_s1;
  --local readdatavalid cpu_data_master_read_data_valid_ddr_sdram_0_s1, which is an e_mux
  cpu_data_master_read_data_valid_ddr_sdram_0_s1 <= ((ddr_sdram_0_s1_readdatavalid_from_sa AND cpu_data_master_rdv_fifo_output_from_ddr_sdram_0_s1)) AND NOT cpu_data_master_rdv_fifo_empty_ddr_sdram_0_s1;
  --ddr_sdram_0_s1_writedata mux, which is an e_mux
  ddr_sdram_0_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ddr_sdram_0_s1)) = '1'), cpu_data_master_writedata, sgdma_rx_m_write_writedata);
  internal_cpu_instruction_master_requests_ddr_sdram_0_s1 <= ((to_std_logic(((Std_Logic_Vector'(cpu_instruction_master_address_to_slave(27 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("0010000000000000000000000000")))) AND (cpu_instruction_master_read))) AND cpu_instruction_master_read;
  --cpu/data_master granted ddr_sdram_0/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_data_master_granted_slave_ddr_sdram_0_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_data_master_granted_slave_ddr_sdram_0_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_data_master_saved_grant_ddr_sdram_0_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((ddr_sdram_0_s1_arbitration_holdoff_internal OR NOT internal_cpu_data_master_requests_ddr_sdram_0_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_data_master_granted_slave_ddr_sdram_0_s1))))));
    end if;

  end process;

  --cpu_data_master_continuerequest continued request, which is an e_mux
  cpu_data_master_continuerequest <= (((last_cycle_cpu_data_master_granted_slave_ddr_sdram_0_s1 AND internal_cpu_data_master_requests_ddr_sdram_0_s1)) OR ((last_cycle_cpu_data_master_granted_slave_ddr_sdram_0_s1 AND internal_cpu_data_master_requests_ddr_sdram_0_s1))) OR ((last_cycle_cpu_data_master_granted_slave_ddr_sdram_0_s1 AND internal_cpu_data_master_requests_ddr_sdram_0_s1));
  internal_cpu_instruction_master_qualified_request_ddr_sdram_0_s1 <= internal_cpu_instruction_master_requests_ddr_sdram_0_s1 AND NOT ((((((cpu_instruction_master_read AND ((to_std_logic(((((std_logic_vector'("00000000000000000000000000000") & (cpu_instruction_master_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("00000000000000000000000000000") & (cpu_instruction_master_latency_counter)))))) OR (cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register))))) OR cpu_data_master_arbiterlock) OR sgdma_rx_m_write_arbiterlock) OR sgdma_tx_m_read_arbiterlock));
  --rdv_fifo_for_cpu_instruction_master_to_ddr_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_ddr_sdram_0_s1 : rdv_fifo_for_cpu_instruction_master_to_ddr_sdram_0_s1_module
    port map(
      data_out => cpu_instruction_master_rdv_fifo_output_from_ddr_sdram_0_s1,
      empty => open,
      fifo_contains_ones_n => cpu_instruction_master_rdv_fifo_empty_ddr_sdram_0_s1,
      full => open,
      clear_fifo => module_input3,
      clk => clk,
      data_in => internal_cpu_instruction_master_granted_ddr_sdram_0_s1,
      read => ddr_sdram_0_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input4,
      write => module_input5
    );

  module_input3 <= std_logic'('0');
  module_input4 <= std_logic'('0');
  module_input5 <= in_a_read_cycle AND NOT ddr_sdram_0_s1_waits_for_read;

  cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register <= NOT cpu_instruction_master_rdv_fifo_empty_ddr_sdram_0_s1;
  --local readdatavalid cpu_instruction_master_read_data_valid_ddr_sdram_0_s1, which is an e_mux
  cpu_instruction_master_read_data_valid_ddr_sdram_0_s1 <= ((ddr_sdram_0_s1_readdatavalid_from_sa AND cpu_instruction_master_rdv_fifo_output_from_ddr_sdram_0_s1)) AND NOT cpu_instruction_master_rdv_fifo_empty_ddr_sdram_0_s1;
  internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_rx_m_write_address_to_slave(31 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000010000000000000000000000000")))) AND (sgdma_rx_m_write_write))) AND sgdma_rx_m_write_write;
  internal_sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 <= internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1 AND NOT (((cpu_data_master_arbiterlock OR cpu_instruction_master_arbiterlock) OR sgdma_tx_m_read_arbiterlock));
  internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_tx_m_read_address_to_slave(31 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("00000010000000000000000000000000")))) AND (sgdma_tx_m_read_read))) AND sgdma_tx_m_read_read;
  internal_sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 <= internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1 AND NOT ((((((sgdma_tx_m_read_read AND to_std_logic((((((std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_m_read_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_m_read_latency_counter))))))))) OR cpu_data_master_arbiterlock) OR cpu_instruction_master_arbiterlock) OR sgdma_rx_m_write_arbiterlock));
  --rdv_fifo_for_sgdma_tx_m_read_to_ddr_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_sgdma_tx_m_read_to_ddr_sdram_0_s1 : rdv_fifo_for_sgdma_tx_m_read_to_ddr_sdram_0_s1_module
    port map(
      data_out => sgdma_tx_m_read_rdv_fifo_output_from_ddr_sdram_0_s1,
      empty => open,
      fifo_contains_ones_n => sgdma_tx_m_read_rdv_fifo_empty_ddr_sdram_0_s1,
      full => open,
      clear_fifo => module_input6,
      clk => clk,
      data_in => internal_sgdma_tx_m_read_granted_ddr_sdram_0_s1,
      read => ddr_sdram_0_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input7,
      write => module_input8
    );

  module_input6 <= std_logic'('0');
  module_input7 <= std_logic'('0');
  module_input8 <= in_a_read_cycle AND NOT ddr_sdram_0_s1_waits_for_read;

  sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register <= NOT sgdma_tx_m_read_rdv_fifo_empty_ddr_sdram_0_s1;
  --local readdatavalid sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1, which is an e_mux
  sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1 <= ((ddr_sdram_0_s1_readdatavalid_from_sa AND sgdma_tx_m_read_rdv_fifo_output_from_ddr_sdram_0_s1)) AND NOT sgdma_tx_m_read_rdv_fifo_empty_ddr_sdram_0_s1;
  --allow new arb cycle for ddr_sdram_0/s1, which is an e_assign
  ddr_sdram_0_s1_allow_new_arb_cycle <= ((NOT cpu_data_master_arbiterlock AND NOT cpu_instruction_master_arbiterlock) AND NOT sgdma_rx_m_write_arbiterlock) AND NOT sgdma_tx_m_read_arbiterlock;
  --sgdma_tx/m_read assignment into master qualified-requests vector for ddr_sdram_0/s1, which is an e_assign
  ddr_sdram_0_s1_master_qreq_vector(0) <= internal_sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1;
  --sgdma_tx/m_read grant ddr_sdram_0/s1, which is an e_assign
  internal_sgdma_tx_m_read_granted_ddr_sdram_0_s1 <= ddr_sdram_0_s1_grant_vector(0);
  --sgdma_tx/m_read saved-grant ddr_sdram_0/s1, which is an e_assign
  sgdma_tx_m_read_saved_grant_ddr_sdram_0_s1 <= ddr_sdram_0_s1_arb_winner(0) AND internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1;
  --sgdma_rx/m_write assignment into master qualified-requests vector for ddr_sdram_0/s1, which is an e_assign
  ddr_sdram_0_s1_master_qreq_vector(1) <= internal_sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1;
  --sgdma_rx/m_write grant ddr_sdram_0/s1, which is an e_assign
  internal_sgdma_rx_m_write_granted_ddr_sdram_0_s1 <= ddr_sdram_0_s1_grant_vector(1);
  --sgdma_rx/m_write saved-grant ddr_sdram_0/s1, which is an e_assign
  sgdma_rx_m_write_saved_grant_ddr_sdram_0_s1 <= ddr_sdram_0_s1_arb_winner(1) AND internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1;
  --cpu/instruction_master assignment into master qualified-requests vector for ddr_sdram_0/s1, which is an e_assign
  ddr_sdram_0_s1_master_qreq_vector(2) <= internal_cpu_instruction_master_qualified_request_ddr_sdram_0_s1;
  --cpu/instruction_master grant ddr_sdram_0/s1, which is an e_assign
  internal_cpu_instruction_master_granted_ddr_sdram_0_s1 <= ddr_sdram_0_s1_grant_vector(2);
  --cpu/instruction_master saved-grant ddr_sdram_0/s1, which is an e_assign
  cpu_instruction_master_saved_grant_ddr_sdram_0_s1 <= ddr_sdram_0_s1_arb_winner(2) AND internal_cpu_instruction_master_requests_ddr_sdram_0_s1;
  --cpu/data_master assignment into master qualified-requests vector for ddr_sdram_0/s1, which is an e_assign
  ddr_sdram_0_s1_master_qreq_vector(3) <= internal_cpu_data_master_qualified_request_ddr_sdram_0_s1;
  --cpu/data_master grant ddr_sdram_0/s1, which is an e_assign
  internal_cpu_data_master_granted_ddr_sdram_0_s1 <= ddr_sdram_0_s1_grant_vector(3);
  --cpu/data_master saved-grant ddr_sdram_0/s1, which is an e_assign
  cpu_data_master_saved_grant_ddr_sdram_0_s1 <= ddr_sdram_0_s1_arb_winner(3) AND internal_cpu_data_master_requests_ddr_sdram_0_s1;
  --ddr_sdram_0/s1 chosen-master double-vector, which is an e_assign
  ddr_sdram_0_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((ddr_sdram_0_s1_master_qreq_vector & ddr_sdram_0_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT ddr_sdram_0_s1_master_qreq_vector & NOT ddr_sdram_0_s1_master_qreq_vector))) + (std_logic_vector'("00000") & (ddr_sdram_0_s1_arb_addend))))), 8);
  --stable onehot encoding of arb winner
  ddr_sdram_0_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((ddr_sdram_0_s1_allow_new_arb_cycle AND or_reduce(ddr_sdram_0_s1_grant_vector)))) = '1'), ddr_sdram_0_s1_grant_vector, ddr_sdram_0_s1_saved_chosen_master_vector);
  --saved ddr_sdram_0_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ddr_sdram_0_s1_saved_chosen_master_vector <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(ddr_sdram_0_s1_allow_new_arb_cycle) = '1' then 
        ddr_sdram_0_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(ddr_sdram_0_s1_grant_vector)) = '1'), ddr_sdram_0_s1_grant_vector, ddr_sdram_0_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  ddr_sdram_0_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((ddr_sdram_0_s1_chosen_master_double_vector(3) OR ddr_sdram_0_s1_chosen_master_double_vector(7)))) & A_ToStdLogicVector(((ddr_sdram_0_s1_chosen_master_double_vector(2) OR ddr_sdram_0_s1_chosen_master_double_vector(6)))) & A_ToStdLogicVector(((ddr_sdram_0_s1_chosen_master_double_vector(1) OR ddr_sdram_0_s1_chosen_master_double_vector(5)))) & A_ToStdLogicVector(((ddr_sdram_0_s1_chosen_master_double_vector(0) OR ddr_sdram_0_s1_chosen_master_double_vector(4)))));
  --ddr_sdram_0/s1 chosen master rotated left, which is an e_assign
  ddr_sdram_0_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(ddr_sdram_0_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("0000")), (std_logic_vector'("0000000000000000000000000000") & ((A_SLL(ddr_sdram_0_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 4);
  --ddr_sdram_0/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ddr_sdram_0_s1_arb_addend <= std_logic_vector'("0001");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(ddr_sdram_0_s1_grant_vector)) = '1' then 
        ddr_sdram_0_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(ddr_sdram_0_s1_end_xfer) = '1'), ddr_sdram_0_s1_chosen_master_rot_left, ddr_sdram_0_s1_grant_vector);
      end if;
    end if;

  end process;

  --ddr_sdram_0_s1_reset_n assignment, which is an e_assign
  ddr_sdram_0_s1_reset_n <= reset_n;
  --ddr_sdram_0_s1_firsttransfer first transaction, which is an e_assign
  ddr_sdram_0_s1_firsttransfer <= A_WE_StdLogic((std_logic'(ddr_sdram_0_s1_begins_xfer) = '1'), ddr_sdram_0_s1_unreg_firsttransfer, ddr_sdram_0_s1_reg_firsttransfer);
  --ddr_sdram_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  ddr_sdram_0_s1_unreg_firsttransfer <= NOT ((ddr_sdram_0_s1_slavearbiterlockenable AND ddr_sdram_0_s1_any_continuerequest));
  --ddr_sdram_0_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ddr_sdram_0_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(ddr_sdram_0_s1_begins_xfer) = '1' then 
        ddr_sdram_0_s1_reg_firsttransfer <= ddr_sdram_0_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --ddr_sdram_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  ddr_sdram_0_s1_beginbursttransfer_internal <= ddr_sdram_0_s1_begins_xfer;
  --ddr_sdram_0_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  ddr_sdram_0_s1_arbitration_holdoff_internal <= ddr_sdram_0_s1_begins_xfer AND ddr_sdram_0_s1_firsttransfer;
  --ddr_sdram_0_s1_read assignment, which is an e_mux
  ddr_sdram_0_s1_read <= (((internal_cpu_data_master_granted_ddr_sdram_0_s1 AND cpu_data_master_read)) OR ((internal_cpu_instruction_master_granted_ddr_sdram_0_s1 AND cpu_instruction_master_read))) OR ((internal_sgdma_tx_m_read_granted_ddr_sdram_0_s1 AND sgdma_tx_m_read_read));
  --ddr_sdram_0_s1_write assignment, which is an e_mux
  ddr_sdram_0_s1_write <= ((internal_cpu_data_master_granted_ddr_sdram_0_s1 AND cpu_data_master_write)) OR ((internal_sgdma_rx_m_write_granted_ddr_sdram_0_s1 AND sgdma_rx_m_write_write));
  shifted_address_to_ddr_sdram_0_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --ddr_sdram_0_s1_address mux, which is an e_mux
  ddr_sdram_0_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ddr_sdram_0_s1)) = '1'), (std_logic_vector'("0000") & ((A_SRL(shifted_address_to_ddr_sdram_0_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010"))))), A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_ddr_sdram_0_s1)) = '1'), (std_logic_vector'("0000") & ((A_SRL(shifted_address_to_ddr_sdram_0_s1_from_cpu_instruction_master,std_logic_vector'("00000000000000000000000000000010"))))), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_m_write_granted_ddr_sdram_0_s1)) = '1'), (A_SRL(shifted_address_to_ddr_sdram_0_s1_from_sgdma_rx_m_write,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_ddr_sdram_0_s1_from_sgdma_tx_m_read,std_logic_vector'("00000000000000000000000000000010")))))), 23);
  shifted_address_to_ddr_sdram_0_s1_from_cpu_instruction_master <= cpu_instruction_master_address_to_slave;
  shifted_address_to_ddr_sdram_0_s1_from_sgdma_rx_m_write <= sgdma_rx_m_write_address_to_slave;
  shifted_address_to_ddr_sdram_0_s1_from_sgdma_tx_m_read <= sgdma_tx_m_read_address_to_slave;
  --d1_ddr_sdram_0_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_ddr_sdram_0_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_ddr_sdram_0_s1_end_xfer <= ddr_sdram_0_s1_end_xfer;
    end if;

  end process;

  --ddr_sdram_0_s1_waits_for_read in a cycle, which is an e_mux
  ddr_sdram_0_s1_waits_for_read <= ddr_sdram_0_s1_in_a_read_cycle AND NOT internal_ddr_sdram_0_s1_waitrequest_n_from_sa;
  --ddr_sdram_0_s1_in_a_read_cycle assignment, which is an e_assign
  ddr_sdram_0_s1_in_a_read_cycle <= (((internal_cpu_data_master_granted_ddr_sdram_0_s1 AND cpu_data_master_read)) OR ((internal_cpu_instruction_master_granted_ddr_sdram_0_s1 AND cpu_instruction_master_read))) OR ((internal_sgdma_tx_m_read_granted_ddr_sdram_0_s1 AND sgdma_tx_m_read_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= ddr_sdram_0_s1_in_a_read_cycle;
  --ddr_sdram_0_s1_waits_for_write in a cycle, which is an e_mux
  ddr_sdram_0_s1_waits_for_write <= ddr_sdram_0_s1_in_a_write_cycle AND NOT internal_ddr_sdram_0_s1_waitrequest_n_from_sa;
  --ddr_sdram_0_s1_in_a_write_cycle assignment, which is an e_assign
  ddr_sdram_0_s1_in_a_write_cycle <= ((internal_cpu_data_master_granted_ddr_sdram_0_s1 AND cpu_data_master_write)) OR ((internal_sgdma_rx_m_write_granted_ddr_sdram_0_s1 AND sgdma_rx_m_write_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= ddr_sdram_0_s1_in_a_write_cycle;
  wait_for_ddr_sdram_0_s1_counter <= std_logic'('0');
  --ddr_sdram_0_s1_byteenable byte enable port mux, which is an e_mux
  ddr_sdram_0_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ddr_sdram_0_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_m_write_granted_ddr_sdram_0_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (sgdma_rx_m_write_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001")))), 4);
  --vhdl renameroo for output signals
  cpu_data_master_granted_ddr_sdram_0_s1 <= internal_cpu_data_master_granted_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_ddr_sdram_0_s1 <= internal_cpu_data_master_qualified_request_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_ddr_sdram_0_s1 <= internal_cpu_data_master_requests_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  cpu_instruction_master_granted_ddr_sdram_0_s1 <= internal_cpu_instruction_master_granted_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  cpu_instruction_master_qualified_request_ddr_sdram_0_s1 <= internal_cpu_instruction_master_qualified_request_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  cpu_instruction_master_requests_ddr_sdram_0_s1 <= internal_cpu_instruction_master_requests_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  ddr_sdram_0_s1_waitrequest_n_from_sa <= internal_ddr_sdram_0_s1_waitrequest_n_from_sa;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_granted_ddr_sdram_0_s1 <= internal_sgdma_rx_m_write_granted_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 <= internal_sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_requests_ddr_sdram_0_s1 <= internal_sgdma_rx_m_write_requests_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_granted_ddr_sdram_0_s1 <= internal_sgdma_tx_m_read_granted_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 <= internal_sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_requests_ddr_sdram_0_s1 <= internal_sgdma_tx_m_read_requests_ddr_sdram_0_s1;
--synthesis translate_off
    --ddr_sdram_0/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line21 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("0000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_data_master_granted_ddr_sdram_0_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_instruction_master_granted_ddr_sdram_0_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(internal_sgdma_rx_m_write_granted_ddr_sdram_0_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_m_read_granted_ddr_sdram_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line21, now);
          write(write_line21, string'(": "));
          write(write_line21, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line21.all);
          deallocate (write_line21);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line22 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("0000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_data_master_saved_grant_ddr_sdram_0_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_saved_grant_ddr_sdram_0_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(sgdma_rx_m_write_saved_grant_ddr_sdram_0_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(sgdma_tx_m_read_saved_grant_ddr_sdram_0_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line22, now);
          write(write_line22, string'(": "));
          write(write_line22, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line22.all);
          deallocate (write_line22);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity descriptor_memory_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_read_latency_counter : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_read : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_write_write : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_read_latency_counter : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_read : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_write_write : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal cpu_data_master_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal d1_descriptor_memory_s1_end_xfer : OUT STD_LOGIC;
                 signal descriptor_memory_s1_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                 signal descriptor_memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal descriptor_memory_s1_chipselect : OUT STD_LOGIC;
                 signal descriptor_memory_s1_clken : OUT STD_LOGIC;
                 signal descriptor_memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal descriptor_memory_s1_write : OUT STD_LOGIC;
                 signal descriptor_memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_read_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_write_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_write_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_write_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_write_requests_descriptor_memory_s1 : OUT STD_LOGIC
              );
end entity descriptor_memory_s1_arbitrator;


architecture europa of descriptor_memory_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in :  STD_LOGIC;
                signal cpu_data_master_saved_grant_descriptor_memory_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal descriptor_memory_s1_allgrants :  STD_LOGIC;
                signal descriptor_memory_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal descriptor_memory_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal descriptor_memory_s1_any_continuerequest :  STD_LOGIC;
                signal descriptor_memory_s1_arb_addend :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_memory_s1_arb_counter_enable :  STD_LOGIC;
                signal descriptor_memory_s1_arb_share_counter :  STD_LOGIC;
                signal descriptor_memory_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal descriptor_memory_s1_arb_share_set_values :  STD_LOGIC;
                signal descriptor_memory_s1_arb_winner :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_memory_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal descriptor_memory_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal descriptor_memory_s1_begins_xfer :  STD_LOGIC;
                signal descriptor_memory_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (9 DOWNTO 0);
                signal descriptor_memory_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_memory_s1_end_xfer :  STD_LOGIC;
                signal descriptor_memory_s1_firsttransfer :  STD_LOGIC;
                signal descriptor_memory_s1_grant_vector :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_memory_s1_in_a_read_cycle :  STD_LOGIC;
                signal descriptor_memory_s1_in_a_write_cycle :  STD_LOGIC;
                signal descriptor_memory_s1_master_qreq_vector :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_memory_s1_non_bursting_master_requests :  STD_LOGIC;
                signal descriptor_memory_s1_reg_firsttransfer :  STD_LOGIC;
                signal descriptor_memory_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal descriptor_memory_s1_slavearbiterlockenable :  STD_LOGIC;
                signal descriptor_memory_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal descriptor_memory_s1_unreg_firsttransfer :  STD_LOGIC;
                signal descriptor_memory_s1_waits_for_read :  STD_LOGIC;
                signal descriptor_memory_s1_waits_for_write :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_descriptor_memory_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_read_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_write_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_read_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_write_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 :  STD_LOGIC;
                signal p1_cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register :  STD_LOGIC;
                signal p1_sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register :  STD_LOGIC;
                signal p1_sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_arbiterlock :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_arbiterlock2 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_continuerequest :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_arbiterlock :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_arbiterlock2 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_continuerequest :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_arbiterlock :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_arbiterlock2 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_continuerequest :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_arbiterlock :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_arbiterlock2 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_continuerequest :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1 :  STD_LOGIC;
                signal shifted_address_to_descriptor_memory_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal wait_for_descriptor_memory_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT descriptor_memory_s1_end_xfer;
    end if;

  end process;

  descriptor_memory_s1_begins_xfer <= NOT d1_reasons_to_wait AND (((((internal_cpu_data_master_qualified_request_descriptor_memory_s1 OR internal_sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1));
  --assign descriptor_memory_s1_readdata_from_sa = descriptor_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  descriptor_memory_s1_readdata_from_sa <= descriptor_memory_s1_readdata;
  internal_cpu_data_master_requests_descriptor_memory_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(27 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("1000010000010000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --descriptor_memory_s1_arb_share_counter set values, which is an e_mux
  descriptor_memory_s1_arb_share_set_values <= std_logic'('1');
  --descriptor_memory_s1_non_bursting_master_requests mux, which is an e_mux
  descriptor_memory_s1_non_bursting_master_requests <= (((((((((((((((((((((((internal_cpu_data_master_requests_descriptor_memory_s1 OR internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1) OR internal_cpu_data_master_requests_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1) OR internal_cpu_data_master_requests_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1) OR internal_cpu_data_master_requests_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1) OR internal_cpu_data_master_requests_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
  --descriptor_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  descriptor_memory_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --descriptor_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  descriptor_memory_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(descriptor_memory_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_memory_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(descriptor_memory_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_memory_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --descriptor_memory_s1_allgrants all slave grants, which is an e_mux
  descriptor_memory_s1_allgrants <= ((((((((((((((((((((((((or_reduce(descriptor_memory_s1_grant_vector)) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector))) OR (or_reduce(descriptor_memory_s1_grant_vector));
  --descriptor_memory_s1_end_xfer assignment, which is an e_assign
  descriptor_memory_s1_end_xfer <= NOT ((descriptor_memory_s1_waits_for_read OR descriptor_memory_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_descriptor_memory_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_descriptor_memory_s1 <= descriptor_memory_s1_end_xfer AND (((NOT descriptor_memory_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --descriptor_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  descriptor_memory_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_descriptor_memory_s1 AND descriptor_memory_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_descriptor_memory_s1 AND NOT descriptor_memory_s1_non_bursting_master_requests));
  --descriptor_memory_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_memory_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(descriptor_memory_s1_arb_counter_enable) = '1' then 
        descriptor_memory_s1_arb_share_counter <= descriptor_memory_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --descriptor_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_memory_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(descriptor_memory_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_descriptor_memory_s1)) OR ((end_xfer_arb_share_counter_term_descriptor_memory_s1 AND NOT descriptor_memory_s1_non_bursting_master_requests)))) = '1' then 
        descriptor_memory_s1_slavearbiterlockenable <= descriptor_memory_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu/data_master descriptor_memory/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= descriptor_memory_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --descriptor_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  descriptor_memory_s1_slavearbiterlockenable2 <= descriptor_memory_s1_arb_share_counter_next_value;
  --cpu/data_master descriptor_memory/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= descriptor_memory_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --sgdma_rx/descriptor_read descriptor_memory/s1 arbiterlock, which is an e_assign
  sgdma_rx_descriptor_read_arbiterlock <= descriptor_memory_s1_slavearbiterlockenable AND sgdma_rx_descriptor_read_continuerequest;
  --sgdma_rx/descriptor_read descriptor_memory/s1 arbiterlock2, which is an e_assign
  sgdma_rx_descriptor_read_arbiterlock2 <= descriptor_memory_s1_slavearbiterlockenable2 AND sgdma_rx_descriptor_read_continuerequest;
  --sgdma_rx/descriptor_read granted descriptor_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_memory_s1_arbitration_holdoff_internal OR NOT internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1))))));
    end if;

  end process;

  --sgdma_rx_descriptor_read_continuerequest continued request, which is an e_mux
  sgdma_rx_descriptor_read_continuerequest <= ((((last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 AND internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1)) OR ((last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 AND internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1))) OR ((last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 AND internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1))) OR ((last_cycle_sgdma_rx_descriptor_read_granted_slave_descriptor_memory_s1 AND internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1));
  --descriptor_memory_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  descriptor_memory_s1_any_continuerequest <= ((((((((((((((((((sgdma_rx_descriptor_read_continuerequest OR sgdma_rx_descriptor_write_continuerequest) OR sgdma_tx_descriptor_read_continuerequest) OR sgdma_tx_descriptor_write_continuerequest) OR cpu_data_master_continuerequest) OR sgdma_rx_descriptor_write_continuerequest) OR sgdma_tx_descriptor_read_continuerequest) OR sgdma_tx_descriptor_write_continuerequest) OR cpu_data_master_continuerequest) OR sgdma_rx_descriptor_read_continuerequest) OR sgdma_tx_descriptor_read_continuerequest) OR sgdma_tx_descriptor_write_continuerequest) OR cpu_data_master_continuerequest) OR sgdma_rx_descriptor_read_continuerequest) OR sgdma_rx_descriptor_write_continuerequest) OR sgdma_tx_descriptor_write_continuerequest) OR cpu_data_master_continuerequest) OR sgdma_rx_descriptor_read_continuerequest) OR sgdma_rx_descriptor_write_continuerequest) OR sgdma_tx_descriptor_read_continuerequest;
  --sgdma_rx/descriptor_write descriptor_memory/s1 arbiterlock, which is an e_assign
  sgdma_rx_descriptor_write_arbiterlock <= descriptor_memory_s1_slavearbiterlockenable AND sgdma_rx_descriptor_write_continuerequest;
  --sgdma_rx/descriptor_write descriptor_memory/s1 arbiterlock2, which is an e_assign
  sgdma_rx_descriptor_write_arbiterlock2 <= descriptor_memory_s1_slavearbiterlockenable2 AND sgdma_rx_descriptor_write_continuerequest;
  --sgdma_rx/descriptor_write granted descriptor_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_memory_s1_arbitration_holdoff_internal OR NOT internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1))))));
    end if;

  end process;

  --sgdma_rx_descriptor_write_continuerequest continued request, which is an e_mux
  sgdma_rx_descriptor_write_continuerequest <= ((((last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 AND internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1)) OR ((last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 AND internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1))) OR ((last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 AND internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1))) OR ((last_cycle_sgdma_rx_descriptor_write_granted_slave_descriptor_memory_s1 AND internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1));
  --sgdma_tx/descriptor_read descriptor_memory/s1 arbiterlock, which is an e_assign
  sgdma_tx_descriptor_read_arbiterlock <= descriptor_memory_s1_slavearbiterlockenable AND sgdma_tx_descriptor_read_continuerequest;
  --sgdma_tx/descriptor_read descriptor_memory/s1 arbiterlock2, which is an e_assign
  sgdma_tx_descriptor_read_arbiterlock2 <= descriptor_memory_s1_slavearbiterlockenable2 AND sgdma_tx_descriptor_read_continuerequest;
  --sgdma_tx/descriptor_read granted descriptor_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_memory_s1_arbitration_holdoff_internal OR NOT internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1))))));
    end if;

  end process;

  --sgdma_tx_descriptor_read_continuerequest continued request, which is an e_mux
  sgdma_tx_descriptor_read_continuerequest <= ((((last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 AND internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1)) OR ((last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 AND internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1))) OR ((last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 AND internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1))) OR ((last_cycle_sgdma_tx_descriptor_read_granted_slave_descriptor_memory_s1 AND internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1));
  --sgdma_tx/descriptor_write descriptor_memory/s1 arbiterlock, which is an e_assign
  sgdma_tx_descriptor_write_arbiterlock <= descriptor_memory_s1_slavearbiterlockenable AND sgdma_tx_descriptor_write_continuerequest;
  --sgdma_tx/descriptor_write descriptor_memory/s1 arbiterlock2, which is an e_assign
  sgdma_tx_descriptor_write_arbiterlock2 <= descriptor_memory_s1_slavearbiterlockenable2 AND sgdma_tx_descriptor_write_continuerequest;
  --sgdma_tx/descriptor_write granted descriptor_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_memory_s1_arbitration_holdoff_internal OR NOT internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1))))));
    end if;

  end process;

  --sgdma_tx_descriptor_write_continuerequest continued request, which is an e_mux
  sgdma_tx_descriptor_write_continuerequest <= ((((last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 AND internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1)) OR ((last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 AND internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1))) OR ((last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 AND internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1))) OR ((last_cycle_sgdma_tx_descriptor_write_granted_slave_descriptor_memory_s1 AND internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1));
  internal_cpu_data_master_qualified_request_descriptor_memory_s1 <= internal_cpu_data_master_requests_descriptor_memory_s1 AND NOT (((((((cpu_data_master_read AND (((to_std_logic(((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("00000000000000000000000000000") & (cpu_data_master_latency_counter))))) OR (cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register)) OR (cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register))))) OR sgdma_rx_descriptor_read_arbiterlock) OR sgdma_rx_descriptor_write_arbiterlock) OR sgdma_tx_descriptor_read_arbiterlock) OR sgdma_tx_descriptor_write_arbiterlock));
  --cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in <= (internal_cpu_data_master_granted_descriptor_memory_s1 AND cpu_data_master_read) AND NOT descriptor_memory_s1_waits_for_read;
  --shift register p1 cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register) & A_ToStdLogicVector(cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register_in)));
  --cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register <= p1_cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_data_master_read_data_valid_descriptor_memory_s1, which is an e_mux
  cpu_data_master_read_data_valid_descriptor_memory_s1 <= cpu_data_master_read_data_valid_descriptor_memory_s1_shift_register;
  --descriptor_memory_s1_writedata mux, which is an e_mux
  descriptor_memory_s1_writedata <= A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_descriptor_memory_s1)) = '1'), cpu_data_master_writedata, A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_write_granted_descriptor_memory_s1)) = '1'), sgdma_rx_descriptor_write_writedata, sgdma_tx_descriptor_write_writedata));
  --mux descriptor_memory_s1_clken, which is an e_mux
  descriptor_memory_s1_clken <= std_logic'('1');
  internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_rx_descriptor_read_address_to_slave(31 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("00001000010000010000000000000000")))) AND (sgdma_rx_descriptor_read_read))) AND sgdma_rx_descriptor_read_read;
  --cpu/data_master granted descriptor_memory/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_data_master_saved_grant_descriptor_memory_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((descriptor_memory_s1_arbitration_holdoff_internal OR NOT internal_cpu_data_master_requests_descriptor_memory_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1))))));
    end if;

  end process;

  --cpu_data_master_continuerequest continued request, which is an e_mux
  cpu_data_master_continuerequest <= ((((last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 AND internal_cpu_data_master_requests_descriptor_memory_s1)) OR ((last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 AND internal_cpu_data_master_requests_descriptor_memory_s1))) OR ((last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 AND internal_cpu_data_master_requests_descriptor_memory_s1))) OR ((last_cycle_cpu_data_master_granted_slave_descriptor_memory_s1 AND internal_cpu_data_master_requests_descriptor_memory_s1));
  internal_sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 <= internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1 AND NOT ((((cpu_data_master_arbiterlock OR sgdma_rx_descriptor_write_arbiterlock) OR sgdma_tx_descriptor_read_arbiterlock) OR sgdma_tx_descriptor_write_arbiterlock));
  --sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in <= (internal_sgdma_rx_descriptor_read_granted_descriptor_memory_s1 AND sgdma_rx_descriptor_read_read) AND NOT descriptor_memory_s1_waits_for_read;
  --shift register p1 sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register) & A_ToStdLogicVector(sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in)));
  --sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= p1_sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1, which is an e_mux
  sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1 <= sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
  internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_rx_descriptor_write_address_to_slave(31 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("00001000010000010000000000000000")))) AND (sgdma_rx_descriptor_write_write))) AND sgdma_rx_descriptor_write_write;
  internal_sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 <= internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1 AND NOT ((((cpu_data_master_arbiterlock OR sgdma_rx_descriptor_read_arbiterlock) OR sgdma_tx_descriptor_read_arbiterlock) OR sgdma_tx_descriptor_write_arbiterlock));
  internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_tx_descriptor_read_address_to_slave(31 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("00001000010000010000000000000000")))) AND (sgdma_tx_descriptor_read_read))) AND sgdma_tx_descriptor_read_read;
  internal_sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 <= internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1 AND NOT ((((cpu_data_master_arbiterlock OR sgdma_rx_descriptor_read_arbiterlock) OR sgdma_rx_descriptor_write_arbiterlock) OR sgdma_tx_descriptor_write_arbiterlock));
  --sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in <= (internal_sgdma_tx_descriptor_read_granted_descriptor_memory_s1 AND sgdma_tx_descriptor_read_read) AND NOT descriptor_memory_s1_waits_for_read;
  --shift register p1 sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register) & A_ToStdLogicVector(sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register_in)));
  --sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register <= p1_sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1, which is an e_mux
  sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1 <= sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1_shift_register;
  internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_tx_descriptor_write_address_to_slave(31 DOWNTO 13) & std_logic_vector'("0000000000000")) = std_logic_vector'("00001000010000010000000000000000")))) AND (sgdma_tx_descriptor_write_write))) AND sgdma_tx_descriptor_write_write;
  internal_sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 <= internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1 AND NOT ((((cpu_data_master_arbiterlock OR sgdma_rx_descriptor_read_arbiterlock) OR sgdma_rx_descriptor_write_arbiterlock) OR sgdma_tx_descriptor_read_arbiterlock));
  --allow new arb cycle for descriptor_memory/s1, which is an e_assign
  descriptor_memory_s1_allow_new_arb_cycle <= (((NOT cpu_data_master_arbiterlock AND NOT sgdma_rx_descriptor_read_arbiterlock) AND NOT sgdma_rx_descriptor_write_arbiterlock) AND NOT sgdma_tx_descriptor_read_arbiterlock) AND NOT sgdma_tx_descriptor_write_arbiterlock;
  --sgdma_tx/descriptor_write assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  descriptor_memory_s1_master_qreq_vector(0) <= internal_sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;
  --sgdma_tx/descriptor_write grant descriptor_memory/s1, which is an e_assign
  internal_sgdma_tx_descriptor_write_granted_descriptor_memory_s1 <= descriptor_memory_s1_grant_vector(0);
  --sgdma_tx/descriptor_write saved-grant descriptor_memory/s1, which is an e_assign
  sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1 <= descriptor_memory_s1_arb_winner(0) AND internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
  --sgdma_tx/descriptor_read assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  descriptor_memory_s1_master_qreq_vector(1) <= internal_sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;
  --sgdma_tx/descriptor_read grant descriptor_memory/s1, which is an e_assign
  internal_sgdma_tx_descriptor_read_granted_descriptor_memory_s1 <= descriptor_memory_s1_grant_vector(1);
  --sgdma_tx/descriptor_read saved-grant descriptor_memory/s1, which is an e_assign
  sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1 <= descriptor_memory_s1_arb_winner(1) AND internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1;
  --sgdma_rx/descriptor_write assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  descriptor_memory_s1_master_qreq_vector(2) <= internal_sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;
  --sgdma_rx/descriptor_write grant descriptor_memory/s1, which is an e_assign
  internal_sgdma_rx_descriptor_write_granted_descriptor_memory_s1 <= descriptor_memory_s1_grant_vector(2);
  --sgdma_rx/descriptor_write saved-grant descriptor_memory/s1, which is an e_assign
  sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1 <= descriptor_memory_s1_arb_winner(2) AND internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1;
  --sgdma_rx/descriptor_read assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  descriptor_memory_s1_master_qreq_vector(3) <= internal_sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;
  --sgdma_rx/descriptor_read grant descriptor_memory/s1, which is an e_assign
  internal_sgdma_rx_descriptor_read_granted_descriptor_memory_s1 <= descriptor_memory_s1_grant_vector(3);
  --sgdma_rx/descriptor_read saved-grant descriptor_memory/s1, which is an e_assign
  sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1 <= descriptor_memory_s1_arb_winner(3) AND internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1;
  --cpu/data_master assignment into master qualified-requests vector for descriptor_memory/s1, which is an e_assign
  descriptor_memory_s1_master_qreq_vector(4) <= internal_cpu_data_master_qualified_request_descriptor_memory_s1;
  --cpu/data_master grant descriptor_memory/s1, which is an e_assign
  internal_cpu_data_master_granted_descriptor_memory_s1 <= descriptor_memory_s1_grant_vector(4);
  --cpu/data_master saved-grant descriptor_memory/s1, which is an e_assign
  cpu_data_master_saved_grant_descriptor_memory_s1 <= descriptor_memory_s1_arb_winner(4) AND internal_cpu_data_master_requests_descriptor_memory_s1;
  --descriptor_memory/s1 chosen-master double-vector, which is an e_assign
  descriptor_memory_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((descriptor_memory_s1_master_qreq_vector & descriptor_memory_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT descriptor_memory_s1_master_qreq_vector & NOT descriptor_memory_s1_master_qreq_vector))) + (std_logic_vector'("000000") & (descriptor_memory_s1_arb_addend))))), 10);
  --stable onehot encoding of arb winner
  descriptor_memory_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((descriptor_memory_s1_allow_new_arb_cycle AND or_reduce(descriptor_memory_s1_grant_vector)))) = '1'), descriptor_memory_s1_grant_vector, descriptor_memory_s1_saved_chosen_master_vector);
  --saved descriptor_memory_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_memory_s1_saved_chosen_master_vector <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      if std_logic'(descriptor_memory_s1_allow_new_arb_cycle) = '1' then 
        descriptor_memory_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(descriptor_memory_s1_grant_vector)) = '1'), descriptor_memory_s1_grant_vector, descriptor_memory_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  descriptor_memory_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((descriptor_memory_s1_chosen_master_double_vector(4) OR descriptor_memory_s1_chosen_master_double_vector(9)))) & A_ToStdLogicVector(((descriptor_memory_s1_chosen_master_double_vector(3) OR descriptor_memory_s1_chosen_master_double_vector(8)))) & A_ToStdLogicVector(((descriptor_memory_s1_chosen_master_double_vector(2) OR descriptor_memory_s1_chosen_master_double_vector(7)))) & A_ToStdLogicVector(((descriptor_memory_s1_chosen_master_double_vector(1) OR descriptor_memory_s1_chosen_master_double_vector(6)))) & A_ToStdLogicVector(((descriptor_memory_s1_chosen_master_double_vector(0) OR descriptor_memory_s1_chosen_master_double_vector(5)))));
  --descriptor_memory/s1 chosen master rotated left, which is an e_assign
  descriptor_memory_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(descriptor_memory_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00000")), (std_logic_vector'("000000000000000000000000000") & ((A_SLL(descriptor_memory_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 5);
  --descriptor_memory/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_memory_s1_arb_addend <= std_logic_vector'("00001");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(descriptor_memory_s1_grant_vector)) = '1' then 
        descriptor_memory_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(descriptor_memory_s1_end_xfer) = '1'), descriptor_memory_s1_chosen_master_rot_left, descriptor_memory_s1_grant_vector);
      end if;
    end if;

  end process;

  descriptor_memory_s1_chipselect <= (((internal_cpu_data_master_granted_descriptor_memory_s1 OR internal_sgdma_rx_descriptor_read_granted_descriptor_memory_s1) OR internal_sgdma_rx_descriptor_write_granted_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_read_granted_descriptor_memory_s1) OR internal_sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  --descriptor_memory_s1_firsttransfer first transaction, which is an e_assign
  descriptor_memory_s1_firsttransfer <= A_WE_StdLogic((std_logic'(descriptor_memory_s1_begins_xfer) = '1'), descriptor_memory_s1_unreg_firsttransfer, descriptor_memory_s1_reg_firsttransfer);
  --descriptor_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  descriptor_memory_s1_unreg_firsttransfer <= NOT ((descriptor_memory_s1_slavearbiterlockenable AND descriptor_memory_s1_any_continuerequest));
  --descriptor_memory_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      descriptor_memory_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(descriptor_memory_s1_begins_xfer) = '1' then 
        descriptor_memory_s1_reg_firsttransfer <= descriptor_memory_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --descriptor_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  descriptor_memory_s1_beginbursttransfer_internal <= descriptor_memory_s1_begins_xfer;
  --descriptor_memory_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  descriptor_memory_s1_arbitration_holdoff_internal <= descriptor_memory_s1_begins_xfer AND descriptor_memory_s1_firsttransfer;
  --descriptor_memory_s1_write assignment, which is an e_mux
  descriptor_memory_s1_write <= (((internal_cpu_data_master_granted_descriptor_memory_s1 AND cpu_data_master_write)) OR ((internal_sgdma_rx_descriptor_write_granted_descriptor_memory_s1 AND sgdma_rx_descriptor_write_write))) OR ((internal_sgdma_tx_descriptor_write_granted_descriptor_memory_s1 AND sgdma_tx_descriptor_write_write));
  shifted_address_to_descriptor_memory_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --descriptor_memory_s1_address mux, which is an e_mux
  descriptor_memory_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_descriptor_memory_s1)) = '1'), (std_logic_vector'("0000") & ((A_SRL(shifted_address_to_descriptor_memory_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010"))))), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_read_granted_descriptor_memory_s1)) = '1'), (A_SRL(shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read,std_logic_vector'("00000000000000000000000000000010"))), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_write_granted_descriptor_memory_s1)) = '1'), (A_SRL(shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write,std_logic_vector'("00000000000000000000000000000010"))), A_WE_StdLogicVector((std_logic'((internal_sgdma_tx_descriptor_read_granted_descriptor_memory_s1)) = '1'), (A_SRL(shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write,std_logic_vector'("00000000000000000000000000000010"))))))), 11);
  shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_read <= sgdma_rx_descriptor_read_address_to_slave;
  shifted_address_to_descriptor_memory_s1_from_sgdma_rx_descriptor_write <= sgdma_rx_descriptor_write_address_to_slave;
  shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_read <= sgdma_tx_descriptor_read_address_to_slave;
  shifted_address_to_descriptor_memory_s1_from_sgdma_tx_descriptor_write <= sgdma_tx_descriptor_write_address_to_slave;
  --d1_descriptor_memory_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_descriptor_memory_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_descriptor_memory_s1_end_xfer <= descriptor_memory_s1_end_xfer;
    end if;

  end process;

  --descriptor_memory_s1_waits_for_read in a cycle, which is an e_mux
  descriptor_memory_s1_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_memory_s1_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --descriptor_memory_s1_in_a_read_cycle assignment, which is an e_assign
  descriptor_memory_s1_in_a_read_cycle <= (((internal_cpu_data_master_granted_descriptor_memory_s1 AND cpu_data_master_read)) OR ((internal_sgdma_rx_descriptor_read_granted_descriptor_memory_s1 AND sgdma_rx_descriptor_read_read))) OR ((internal_sgdma_tx_descriptor_read_granted_descriptor_memory_s1 AND sgdma_tx_descriptor_read_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= descriptor_memory_s1_in_a_read_cycle;
  --descriptor_memory_s1_waits_for_write in a cycle, which is an e_mux
  descriptor_memory_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(descriptor_memory_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --descriptor_memory_s1_in_a_write_cycle assignment, which is an e_assign
  descriptor_memory_s1_in_a_write_cycle <= (((internal_cpu_data_master_granted_descriptor_memory_s1 AND cpu_data_master_write)) OR ((internal_sgdma_rx_descriptor_write_granted_descriptor_memory_s1 AND sgdma_rx_descriptor_write_write))) OR ((internal_sgdma_tx_descriptor_write_granted_descriptor_memory_s1 AND sgdma_tx_descriptor_write_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= descriptor_memory_s1_in_a_write_cycle;
  wait_for_descriptor_memory_s1_counter <= std_logic'('0');
  --descriptor_memory_s1_byteenable byte enable port mux, which is an e_mux
  descriptor_memory_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_descriptor_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_write_granted_descriptor_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (A_REP(std_logic'('1'), 4))), A_WE_StdLogicVector((std_logic'((internal_sgdma_tx_descriptor_write_granted_descriptor_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (A_REP(std_logic'('1'), 4))), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))))), 4);
  --vhdl renameroo for output signals
  cpu_data_master_granted_descriptor_memory_s1 <= internal_cpu_data_master_granted_descriptor_memory_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_descriptor_memory_s1 <= internal_cpu_data_master_qualified_request_descriptor_memory_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_descriptor_memory_s1 <= internal_cpu_data_master_requests_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_granted_descriptor_memory_s1 <= internal_sgdma_rx_descriptor_read_granted_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 <= internal_sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_requests_descriptor_memory_s1 <= internal_sgdma_rx_descriptor_read_requests_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_write_granted_descriptor_memory_s1 <= internal_sgdma_rx_descriptor_write_granted_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 <= internal_sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_write_requests_descriptor_memory_s1 <= internal_sgdma_rx_descriptor_write_requests_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_granted_descriptor_memory_s1 <= internal_sgdma_tx_descriptor_read_granted_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 <= internal_sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_requests_descriptor_memory_s1 <= internal_sgdma_tx_descriptor_read_requests_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_write_granted_descriptor_memory_s1 <= internal_sgdma_tx_descriptor_write_granted_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 <= internal_sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_write_requests_descriptor_memory_s1 <= internal_sgdma_tx_descriptor_write_requests_descriptor_memory_s1;
--synthesis translate_off
    --descriptor_memory/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line23 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_data_master_granted_descriptor_memory_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_sgdma_rx_descriptor_read_granted_descriptor_memory_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(internal_sgdma_rx_descriptor_write_granted_descriptor_memory_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_descriptor_read_granted_descriptor_memory_s1)))))) + (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_descriptor_write_granted_descriptor_memory_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line23, now);
          write(write_line23, string'(": "));
          write(write_line23, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line23.all);
          deallocate (write_line23);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line24 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_data_master_saved_grant_descriptor_memory_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(sgdma_rx_descriptor_read_saved_grant_descriptor_memory_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(sgdma_rx_descriptor_write_saved_grant_descriptor_memory_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(sgdma_tx_descriptor_read_saved_grant_descriptor_memory_s1)))))) + (std_logic_vector'("0000") & (A_TOSTDLOGICVECTOR(sgdma_tx_descriptor_write_saved_grant_descriptor_memory_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line24, now);
          write(write_line24, string'(": "));
          write(write_line24, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line24.all);
          deallocate (write_line24);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ext_flash_enet_bus_avalon_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_ext_flash_enet_bus_avalon_slave_end_xfer : OUT STD_LOGIC;
                 signal ext_flash_enet_bus_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal ext_flash_enet_bus_data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal ext_flash_s1_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pipeline_bridge_m1_byteenable_ext_flash_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_ext_flash_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_ext_flash_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_ext_flash_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_ext_flash_s1 : OUT STD_LOGIC;
                 signal read_n_to_the_ext_flash : OUT STD_LOGIC;
                 signal select_n_to_the_ext_flash : OUT STD_LOGIC;
                 signal write_n_to_the_ext_flash : OUT STD_LOGIC
              );
end entity ext_flash_enet_bus_avalon_slave_arbitrator;


architecture europa of ext_flash_enet_bus_avalon_slave_arbitrator is
                signal d1_in_a_write_cycle :  STD_LOGIC;
                signal d1_outgoing_ext_flash_enet_bus_data :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_ext_flash_enet_bus_avalon_slave :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_allgrants :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_any_continuerequest :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_arb_counter_enable :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal ext_flash_enet_bus_avalon_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal ext_flash_enet_bus_avalon_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal ext_flash_enet_bus_avalon_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_begins_xfer :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_end_xfer :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_firsttransfer :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_grant_vector :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_master_qreq_vector :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_non_bursting_master_requests :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_read_pending :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_reg_firsttransfer :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_slavearbiterlockenable :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_unreg_firsttransfer :  STD_LOGIC;
                signal ext_flash_enet_bus_avalon_slave_write_pending :  STD_LOGIC;
                signal ext_flash_s1_counter_load_value :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal ext_flash_s1_in_a_read_cycle :  STD_LOGIC;
                signal ext_flash_s1_in_a_write_cycle :  STD_LOGIC;
                signal ext_flash_s1_pretend_byte_enable :  STD_LOGIC;
                signal ext_flash_s1_wait_counter :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal ext_flash_s1_waits_for_read :  STD_LOGIC;
                signal ext_flash_s1_waits_for_write :  STD_LOGIC;
                signal ext_flash_s1_with_write_latency :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal incoming_ext_flash_enet_bus_data :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal incoming_ext_flash_enet_bus_data_bit_0_is_x :  STD_LOGIC;
                signal incoming_ext_flash_enet_bus_data_bit_1_is_x :  STD_LOGIC;
                signal incoming_ext_flash_enet_bus_data_bit_2_is_x :  STD_LOGIC;
                signal incoming_ext_flash_enet_bus_data_bit_3_is_x :  STD_LOGIC;
                signal incoming_ext_flash_enet_bus_data_bit_4_is_x :  STD_LOGIC;
                signal incoming_ext_flash_enet_bus_data_bit_5_is_x :  STD_LOGIC;
                signal incoming_ext_flash_enet_bus_data_bit_6_is_x :  STD_LOGIC;
                signal incoming_ext_flash_enet_bus_data_bit_7_is_x :  STD_LOGIC;
                signal internal_ext_flash_s1_wait_counter_eq_0 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_byteenable_ext_flash_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_ext_flash_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_ext_flash_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_ext_flash_s1 :  STD_LOGIC;
                signal outgoing_ext_flash_enet_bus_data :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_ext_flash_enet_bus_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal p1_pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_read_n_to_the_ext_flash :  STD_LOGIC;
                signal p1_select_n_to_the_ext_flash :  STD_LOGIC;
                signal p1_write_n_to_the_ext_flash :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_byteenable_ext_flash_s1_segment_0 :  STD_LOGIC;
                signal pipeline_bridge_m1_byteenable_ext_flash_s1_segment_1 :  STD_LOGIC;
                signal pipeline_bridge_m1_byteenable_ext_flash_s1_segment_2 :  STD_LOGIC;
                signal pipeline_bridge_m1_byteenable_ext_flash_s1_segment_3 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register_in :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_ext_flash_s1 :  STD_LOGIC;
                signal time_to_write :  STD_LOGIC;
                signal wait_for_ext_flash_s1_counter :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of d1_in_a_write_cycle : signal is "FAST_OUTPUT_ENABLE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of d1_outgoing_ext_flash_enet_bus_data : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of ext_flash_enet_bus_address : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of incoming_ext_flash_enet_bus_data : signal is "FAST_INPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of read_n_to_the_ext_flash : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of select_n_to_the_ext_flash : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of write_n_to_the_ext_flash : signal is "FAST_OUTPUT_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT ext_flash_enet_bus_avalon_slave_end_xfer;
    end if;

  end process;

  ext_flash_enet_bus_avalon_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_ext_flash_s1);
  internal_pipeline_bridge_m1_requests_ext_flash_s1 <= to_std_logic(((Std_Logic_Vector'(A_ToStdLogicVector(pipeline_bridge_m1_address_to_slave(24)) & std_logic_vector'("000000000000000000000000")) = std_logic_vector'("0000000000000000000000000")))) AND pipeline_bridge_m1_chipselect;
  --~select_n_to_the_ext_flash of type chipselect to ~p1_select_n_to_the_ext_flash, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      select_n_to_the_ext_flash <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      select_n_to_the_ext_flash <= p1_select_n_to_the_ext_flash;
    end if;

  end process;

  ext_flash_enet_bus_avalon_slave_write_pending <= std_logic'('0');
  --ext_flash_enet_bus/avalon_slave read pending calc, which is an e_assign
  ext_flash_enet_bus_avalon_slave_read_pending <= std_logic'('0');
  --ext_flash_enet_bus_avalon_slave_arb_share_counter set values, which is an e_mux
  ext_flash_enet_bus_avalon_slave_arb_share_set_values <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_m1_granted_ext_flash_s1)) = '1'), std_logic_vector'("00000000000000000000000000000100"), std_logic_vector'("00000000000000000000000000000001")), 3);
  --ext_flash_enet_bus_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  ext_flash_enet_bus_avalon_slave_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_ext_flash_s1;
  --ext_flash_enet_bus_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  ext_flash_enet_bus_avalon_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --ext_flash_enet_bus_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  ext_flash_enet_bus_avalon_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(ext_flash_enet_bus_avalon_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (ext_flash_enet_bus_avalon_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(ext_flash_enet_bus_avalon_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (ext_flash_enet_bus_avalon_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --ext_flash_enet_bus_avalon_slave_allgrants all slave grants, which is an e_mux
  ext_flash_enet_bus_avalon_slave_allgrants <= ext_flash_enet_bus_avalon_slave_grant_vector;
  --ext_flash_enet_bus_avalon_slave_end_xfer assignment, which is an e_assign
  ext_flash_enet_bus_avalon_slave_end_xfer <= NOT ((ext_flash_s1_waits_for_read OR ext_flash_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_ext_flash_enet_bus_avalon_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_ext_flash_enet_bus_avalon_slave <= ext_flash_enet_bus_avalon_slave_end_xfer AND (((NOT ext_flash_enet_bus_avalon_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --ext_flash_enet_bus_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  ext_flash_enet_bus_avalon_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_ext_flash_enet_bus_avalon_slave AND ext_flash_enet_bus_avalon_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_ext_flash_enet_bus_avalon_slave AND NOT ext_flash_enet_bus_avalon_slave_non_bursting_master_requests));
  --ext_flash_enet_bus_avalon_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_flash_enet_bus_avalon_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(ext_flash_enet_bus_avalon_slave_arb_counter_enable) = '1' then 
        ext_flash_enet_bus_avalon_slave_arb_share_counter <= ext_flash_enet_bus_avalon_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ext_flash_enet_bus_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_flash_enet_bus_avalon_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((ext_flash_enet_bus_avalon_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_ext_flash_enet_bus_avalon_slave)) OR ((end_xfer_arb_share_counter_term_ext_flash_enet_bus_avalon_slave AND NOT ext_flash_enet_bus_avalon_slave_non_bursting_master_requests)))) = '1' then 
        ext_flash_enet_bus_avalon_slave_slavearbiterlockenable <= or_reduce(ext_flash_enet_bus_avalon_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 ext_flash_enet_bus/avalon_slave arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= ext_flash_enet_bus_avalon_slave_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --ext_flash_enet_bus_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  ext_flash_enet_bus_avalon_slave_slavearbiterlockenable2 <= or_reduce(ext_flash_enet_bus_avalon_slave_arb_share_counter_next_value);
  --pipeline_bridge/m1 ext_flash_enet_bus/avalon_slave arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= ext_flash_enet_bus_avalon_slave_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --ext_flash_enet_bus_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  ext_flash_enet_bus_avalon_slave_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_ext_flash_s1 <= internal_pipeline_bridge_m1_requests_ext_flash_s1 AND NOT ((((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND (((ext_flash_enet_bus_avalon_slave_write_pending OR (ext_flash_enet_bus_avalon_slave_read_pending)) OR to_std_logic(((std_logic_vector'("00000000000000000000000000000010")<(std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter))))))))) OR ((((ext_flash_enet_bus_avalon_slave_read_pending OR NOT(internal_pipeline_bridge_m1_byteenable_ext_flash_s1))) AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect))))));
  --pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register_in <= (internal_pipeline_bridge_m1_granted_ext_flash_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT ext_flash_s1_waits_for_read;
  --shift register p1 pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register <= A_EXT ((pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register & A_ToStdLogicVector(pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register_in)), 2);
  --pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register <= p1_pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register;
    end if;

  end process;

  --local readdatavalid pipeline_bridge_m1_read_data_valid_ext_flash_s1, which is an e_mux
  pipeline_bridge_m1_read_data_valid_ext_flash_s1 <= pipeline_bridge_m1_read_data_valid_ext_flash_s1_shift_register(1);
  --ext_flash_enet_bus_data register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      incoming_ext_flash_enet_bus_data <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      incoming_ext_flash_enet_bus_data <= ext_flash_enet_bus_data;
    end if;

  end process;

  --ext_flash_s1_with_write_latency assignment, which is an e_assign
  ext_flash_s1_with_write_latency <= in_a_write_cycle AND (internal_pipeline_bridge_m1_qualified_request_ext_flash_s1);
  --time to write the data, which is an e_mux
  time_to_write <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((ext_flash_s1_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), std_logic_vector'("00000000000000000000000000000000")));
  --d1_outgoing_ext_flash_enet_bus_data register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_outgoing_ext_flash_enet_bus_data <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      d1_outgoing_ext_flash_enet_bus_data <= outgoing_ext_flash_enet_bus_data;
    end if;

  end process;

  --write cycle delayed by 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_in_a_write_cycle <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_in_a_write_cycle <= time_to_write;
    end if;

  end process;

  --d1_outgoing_ext_flash_enet_bus_data tristate driver, which is an e_assign
  ext_flash_enet_bus_data <= A_WE_StdLogicVector((std_logic'((d1_in_a_write_cycle)) = '1'), d1_outgoing_ext_flash_enet_bus_data, A_REP(std_logic'('Z'), 8));
  --outgoing_ext_flash_enet_bus_data mux, which is an e_mux
  outgoing_ext_flash_enet_bus_data <= pipeline_bridge_m1_dbs_write_8;
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_ext_flash_s1 <= internal_pipeline_bridge_m1_qualified_request_ext_flash_s1;
  --pipeline_bridge/m1 saved-grant ext_flash/s1, which is an e_assign
  pipeline_bridge_m1_saved_grant_ext_flash_s1 <= internal_pipeline_bridge_m1_requests_ext_flash_s1;
  --allow new arb cycle for ext_flash_enet_bus/avalon_slave, which is an e_assign
  ext_flash_enet_bus_avalon_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  ext_flash_enet_bus_avalon_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  ext_flash_enet_bus_avalon_slave_master_qreq_vector <= std_logic'('1');
  p1_select_n_to_the_ext_flash <= NOT internal_pipeline_bridge_m1_granted_ext_flash_s1;
  --ext_flash_enet_bus_avalon_slave_firsttransfer first transaction, which is an e_assign
  ext_flash_enet_bus_avalon_slave_firsttransfer <= A_WE_StdLogic((std_logic'(ext_flash_enet_bus_avalon_slave_begins_xfer) = '1'), ext_flash_enet_bus_avalon_slave_unreg_firsttransfer, ext_flash_enet_bus_avalon_slave_reg_firsttransfer);
  --ext_flash_enet_bus_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  ext_flash_enet_bus_avalon_slave_unreg_firsttransfer <= NOT ((ext_flash_enet_bus_avalon_slave_slavearbiterlockenable AND ext_flash_enet_bus_avalon_slave_any_continuerequest));
  --ext_flash_enet_bus_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_flash_enet_bus_avalon_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(ext_flash_enet_bus_avalon_slave_begins_xfer) = '1' then 
        ext_flash_enet_bus_avalon_slave_reg_firsttransfer <= ext_flash_enet_bus_avalon_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --ext_flash_enet_bus_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  ext_flash_enet_bus_avalon_slave_beginbursttransfer_internal <= ext_flash_enet_bus_avalon_slave_begins_xfer;
  --~read_n_to_the_ext_flash of type read to ~p1_read_n_to_the_ext_flash, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      read_n_to_the_ext_flash <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      read_n_to_the_ext_flash <= p1_read_n_to_the_ext_flash;
    end if;

  end process;

  --~p1_read_n_to_the_ext_flash assignment, which is an e_mux
  p1_read_n_to_the_ext_flash <= NOT (((((internal_pipeline_bridge_m1_granted_ext_flash_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) AND NOT ext_flash_enet_bus_avalon_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("00000000000000000000000000") & (ext_flash_s1_wait_counter))<std_logic_vector'("00000000000000000000000000011000"))))));
  --~write_n_to_the_ext_flash of type write to ~p1_write_n_to_the_ext_flash, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      write_n_to_the_ext_flash <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      write_n_to_the_ext_flash <= p1_write_n_to_the_ext_flash;
    end if;

  end process;

  --~p1_write_n_to_the_ext_flash assignment, which is an e_mux
  p1_write_n_to_the_ext_flash <= NOT (((((((internal_pipeline_bridge_m1_granted_ext_flash_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))) AND NOT ext_flash_enet_bus_avalon_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("00000000000000000000000000") & (ext_flash_s1_wait_counter))>=std_logic_vector'("00000000000000000000000000000110"))))) AND to_std_logic((((std_logic_vector'("00000000000000000000000000") & (ext_flash_s1_wait_counter))<std_logic_vector'("00000000000000000000000000011110"))))) AND ext_flash_s1_pretend_byte_enable));
  --ext_flash_enet_bus_address of type address to p1_ext_flash_enet_bus_address, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_flash_enet_bus_address <= std_logic_vector'("000000000000000000000000");
    elsif clk'event and clk = '1' then
      ext_flash_enet_bus_address <= p1_ext_flash_enet_bus_address;
    end if;

  end process;

  --p1_ext_flash_enet_bus_address mux, which is an e_mux
  p1_ext_flash_enet_bus_address <= A_EXT (Std_Logic_Vector'(A_SRL(pipeline_bridge_m1_address_to_slave,std_logic_vector'("00000000000000000000000000000010")) & pipeline_bridge_m1_dbs_address(1 DOWNTO 0)), 24);
  --d1_ext_flash_enet_bus_avalon_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_ext_flash_enet_bus_avalon_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_ext_flash_enet_bus_avalon_slave_end_xfer <= ext_flash_enet_bus_avalon_slave_end_xfer;
    end if;

  end process;

  --ext_flash_s1_waits_for_read in a cycle, which is an e_mux
  ext_flash_s1_waits_for_read <= ext_flash_s1_in_a_read_cycle AND wait_for_ext_flash_s1_counter;
  --ext_flash_s1_in_a_read_cycle assignment, which is an e_assign
  ext_flash_s1_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_ext_flash_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= ext_flash_s1_in_a_read_cycle;
  --ext_flash_s1_waits_for_write in a cycle, which is an e_mux
  ext_flash_s1_waits_for_write <= ext_flash_s1_in_a_write_cycle AND wait_for_ext_flash_s1_counter;
  --ext_flash_s1_in_a_write_cycle assignment, which is an e_assign
  ext_flash_s1_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_ext_flash_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= ext_flash_s1_in_a_write_cycle;
  internal_ext_flash_s1_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("00000000000000000000000000") & (ext_flash_s1_wait_counter)) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_flash_s1_wait_counter <= std_logic_vector'("000000");
    elsif clk'event and clk = '1' then
      ext_flash_s1_wait_counter <= ext_flash_s1_counter_load_value;
    end if;

  end process;

  ext_flash_s1_counter_load_value <= A_EXT (A_WE_StdLogicVector((std_logic'(((ext_flash_s1_in_a_read_cycle AND ext_flash_enet_bus_avalon_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000011101"), A_WE_StdLogicVector((std_logic'(((ext_flash_s1_in_a_write_cycle AND ext_flash_enet_bus_avalon_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000000100011"), A_WE_StdLogicVector((std_logic'((NOT internal_ext_flash_s1_wait_counter_eq_0)) = '1'), ((std_logic_vector'("000000000000000000000000000") & (ext_flash_s1_wait_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000")))), 6);
  wait_for_ext_flash_s1_counter <= ext_flash_enet_bus_avalon_slave_begins_xfer OR NOT internal_ext_flash_s1_wait_counter_eq_0;
  --ext_flash_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  ext_flash_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_m1_granted_ext_flash_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_pipeline_bridge_m1_byteenable_ext_flash_s1))), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  (pipeline_bridge_m1_byteenable_ext_flash_s1_segment_3, pipeline_bridge_m1_byteenable_ext_flash_s1_segment_2, pipeline_bridge_m1_byteenable_ext_flash_s1_segment_1, pipeline_bridge_m1_byteenable_ext_flash_s1_segment_0) <= pipeline_bridge_m1_byteenable;
  internal_pipeline_bridge_m1_byteenable_ext_flash_s1 <= A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), pipeline_bridge_m1_byteenable_ext_flash_s1_segment_0, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), pipeline_bridge_m1_byteenable_ext_flash_s1_segment_1, A_WE_StdLogic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), pipeline_bridge_m1_byteenable_ext_flash_s1_segment_2, pipeline_bridge_m1_byteenable_ext_flash_s1_segment_3)));
  --vhdl renameroo for output signals
  ext_flash_s1_wait_counter_eq_0 <= internal_ext_flash_s1_wait_counter_eq_0;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_byteenable_ext_flash_s1 <= internal_pipeline_bridge_m1_byteenable_ext_flash_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_ext_flash_s1 <= internal_pipeline_bridge_m1_granted_ext_flash_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_ext_flash_s1 <= internal_pipeline_bridge_m1_qualified_request_ext_flash_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_ext_flash_s1 <= internal_pipeline_bridge_m1_requests_ext_flash_s1;
--synthesis translate_off
    --incoming_ext_flash_enet_bus_data_bit_0_is_x x check, which is an e_assign_is_x
    incoming_ext_flash_enet_bus_data_bit_0_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_ext_flash_enet_bus_data(0))), '1','0');
    --Crush incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0[0] Xs to 0, which is an e_assign
    incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0(0) <= A_WE_StdLogic((std_logic'(incoming_ext_flash_enet_bus_data_bit_0_is_x) = '1'), std_logic'('0'), incoming_ext_flash_enet_bus_data(0));
    --incoming_ext_flash_enet_bus_data_bit_1_is_x x check, which is an e_assign_is_x
    incoming_ext_flash_enet_bus_data_bit_1_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_ext_flash_enet_bus_data(1))), '1','0');
    --Crush incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0[1] Xs to 0, which is an e_assign
    incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0(1) <= A_WE_StdLogic((std_logic'(incoming_ext_flash_enet_bus_data_bit_1_is_x) = '1'), std_logic'('0'), incoming_ext_flash_enet_bus_data(1));
    --incoming_ext_flash_enet_bus_data_bit_2_is_x x check, which is an e_assign_is_x
    incoming_ext_flash_enet_bus_data_bit_2_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_ext_flash_enet_bus_data(2))), '1','0');
    --Crush incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0[2] Xs to 0, which is an e_assign
    incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0(2) <= A_WE_StdLogic((std_logic'(incoming_ext_flash_enet_bus_data_bit_2_is_x) = '1'), std_logic'('0'), incoming_ext_flash_enet_bus_data(2));
    --incoming_ext_flash_enet_bus_data_bit_3_is_x x check, which is an e_assign_is_x
    incoming_ext_flash_enet_bus_data_bit_3_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_ext_flash_enet_bus_data(3))), '1','0');
    --Crush incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0[3] Xs to 0, which is an e_assign
    incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0(3) <= A_WE_StdLogic((std_logic'(incoming_ext_flash_enet_bus_data_bit_3_is_x) = '1'), std_logic'('0'), incoming_ext_flash_enet_bus_data(3));
    --incoming_ext_flash_enet_bus_data_bit_4_is_x x check, which is an e_assign_is_x
    incoming_ext_flash_enet_bus_data_bit_4_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_ext_flash_enet_bus_data(4))), '1','0');
    --Crush incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0[4] Xs to 0, which is an e_assign
    incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0(4) <= A_WE_StdLogic((std_logic'(incoming_ext_flash_enet_bus_data_bit_4_is_x) = '1'), std_logic'('0'), incoming_ext_flash_enet_bus_data(4));
    --incoming_ext_flash_enet_bus_data_bit_5_is_x x check, which is an e_assign_is_x
    incoming_ext_flash_enet_bus_data_bit_5_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_ext_flash_enet_bus_data(5))), '1','0');
    --Crush incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0[5] Xs to 0, which is an e_assign
    incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0(5) <= A_WE_StdLogic((std_logic'(incoming_ext_flash_enet_bus_data_bit_5_is_x) = '1'), std_logic'('0'), incoming_ext_flash_enet_bus_data(5));
    --incoming_ext_flash_enet_bus_data_bit_6_is_x x check, which is an e_assign_is_x
    incoming_ext_flash_enet_bus_data_bit_6_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_ext_flash_enet_bus_data(6))), '1','0');
    --Crush incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0[6] Xs to 0, which is an e_assign
    incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0(6) <= A_WE_StdLogic((std_logic'(incoming_ext_flash_enet_bus_data_bit_6_is_x) = '1'), std_logic'('0'), incoming_ext_flash_enet_bus_data(6));
    --incoming_ext_flash_enet_bus_data_bit_7_is_x x check, which is an e_assign_is_x
    incoming_ext_flash_enet_bus_data_bit_7_is_x <= A_WE_StdLogic(is_x(std_ulogic(incoming_ext_flash_enet_bus_data(7))), '1','0');
    --Crush incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0[7] Xs to 0, which is an e_assign
    incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0(7) <= A_WE_StdLogic((std_logic'(incoming_ext_flash_enet_bus_data_bit_7_is_x) = '1'), std_logic'('0'), incoming_ext_flash_enet_bus_data(7));
    --ext_flash/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line25 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_ext_flash_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line25, now);
          write(write_line25, string'(": "));
          write(write_line25, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave ext_flash/s1"));
          write(output, write_line25.all);
          deallocate (write_line25);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on
--synthesis read_comments_as_HDL on
--    
--    incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0 <= incoming_ext_flash_enet_bus_data;
--synthesis read_comments_as_HDL off

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ext_flash_enet_bus_bridge_arbitrator is 
end entity ext_flash_enet_bus_bridge_arbitrator;


architecture europa of ext_flash_enet_bus_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ext_ssram_bus_avalon_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_m_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal sgdma_rx_m_write_write : IN STD_LOGIC;
                 signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal sgdma_tx_m_read_read : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;

              -- outputs:
                 signal adsc_n_to_the_ext_ssram : OUT STD_LOGIC;
                 signal bw_n_to_the_ext_ssram : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal bwe_n_to_the_ext_ssram : OUT STD_LOGIC;
                 signal chipenable1_n_to_the_ext_ssram : OUT STD_LOGIC;
                 signal cpu_data_master_granted_ext_ssram_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_ext_ssram_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ext_ssram_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_ext_ssram_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_granted_ext_ssram_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_ext_ssram_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_ext_ssram_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_requests_ext_ssram_s1 : OUT STD_LOGIC;
                 signal d1_ext_ssram_bus_avalon_slave_end_xfer : OUT STD_LOGIC;
                 signal ext_ssram_bus_address : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal ext_ssram_bus_data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal incoming_ext_ssram_bus_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal outputenable_n_to_the_ext_ssram : OUT STD_LOGIC;
                 signal sgdma_rx_m_write_granted_ext_ssram_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_m_write_qualified_request_ext_ssram_s1 : OUT STD_LOGIC;
                 signal sgdma_rx_m_write_requests_ext_ssram_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_granted_ext_ssram_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_qualified_request_ext_ssram_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_ext_ssram_s1 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_requests_ext_ssram_s1 : OUT STD_LOGIC
              );
end entity ext_ssram_bus_avalon_slave_arbitrator;


architecture europa of ext_ssram_bus_avalon_slave_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_ext_ssram_s1_shift_register :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_data_master_read_data_valid_ext_ssram_s1_shift_register_in :  STD_LOGIC;
                signal cpu_data_master_saved_grant_ext_ssram_s1 :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register_in :  STD_LOGIC;
                signal cpu_instruction_master_saved_grant_ext_ssram_s1 :  STD_LOGIC;
                signal d1_in_a_write_cycle :  STD_LOGIC;
                signal d1_outgoing_ext_ssram_bus_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_allgrants :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_any_continuerequest :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_arb_addend :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ext_ssram_bus_avalon_slave_arb_counter_enable :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_arb_share_counter :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_arb_share_counter_next_value :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_arb_share_set_values :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_arb_winner :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ext_ssram_bus_avalon_slave_arbitration_holdoff_internal :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_begins_xfer :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_chosen_master_double_vector :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal ext_ssram_bus_avalon_slave_chosen_master_rot_left :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ext_ssram_bus_avalon_slave_end_xfer :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_firsttransfer :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_grant_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ext_ssram_bus_avalon_slave_master_qreq_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ext_ssram_bus_avalon_slave_non_bursting_master_requests :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_read_pending :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_reg_firsttransfer :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_saved_chosen_master_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ext_ssram_bus_avalon_slave_slavearbiterlockenable :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_unreg_firsttransfer :  STD_LOGIC;
                signal ext_ssram_bus_avalon_slave_write_pending :  STD_LOGIC;
                signal ext_ssram_s1_in_a_read_cycle :  STD_LOGIC;
                signal ext_ssram_s1_in_a_write_cycle :  STD_LOGIC;
                signal ext_ssram_s1_waits_for_read :  STD_LOGIC;
                signal ext_ssram_s1_waits_for_write :  STD_LOGIC;
                signal ext_ssram_s1_with_write_latency :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_ext_ssram_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_ext_ssram_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_ext_ssram_s1 :  STD_LOGIC;
                signal internal_cpu_instruction_master_granted_ext_ssram_s1 :  STD_LOGIC;
                signal internal_cpu_instruction_master_qualified_request_ext_ssram_s1 :  STD_LOGIC;
                signal internal_cpu_instruction_master_requests_ext_ssram_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_granted_ext_ssram_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_qualified_request_ext_ssram_s1 :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_requests_ext_ssram_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_granted_ext_ssram_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_qualified_request_ext_ssram_s1 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_requests_ext_ssram_s1 :  STD_LOGIC;
                signal last_cycle_cpu_data_master_granted_slave_ext_ssram_s1 :  STD_LOGIC;
                signal last_cycle_cpu_instruction_master_granted_slave_ext_ssram_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_rx_m_write_granted_slave_ext_ssram_s1 :  STD_LOGIC;
                signal last_cycle_sgdma_tx_m_read_granted_slave_ext_ssram_s1 :  STD_LOGIC;
                signal outgoing_ext_ssram_bus_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal p1_adsc_n_to_the_ext_ssram :  STD_LOGIC;
                signal p1_bw_n_to_the_ext_ssram :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p1_bwe_n_to_the_ext_ssram :  STD_LOGIC;
                signal p1_chipenable1_n_to_the_ext_ssram :  STD_LOGIC;
                signal p1_cpu_data_master_read_data_valid_ext_ssram_s1_shift_register :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p1_cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal p1_ext_ssram_bus_address :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal p1_outputenable_n_to_the_ext_ssram :  STD_LOGIC;
                signal p1_sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sgdma_rx_m_write_arbiterlock :  STD_LOGIC;
                signal sgdma_rx_m_write_arbiterlock2 :  STD_LOGIC;
                signal sgdma_rx_m_write_continuerequest :  STD_LOGIC;
                signal sgdma_rx_m_write_saved_grant_ext_ssram_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_arbiterlock :  STD_LOGIC;
                signal sgdma_tx_m_read_arbiterlock2 :  STD_LOGIC;
                signal sgdma_tx_m_read_continuerequest :  STD_LOGIC;
                signal sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register_in :  STD_LOGIC;
                signal sgdma_tx_m_read_saved_grant_ext_ssram_s1 :  STD_LOGIC;
                signal time_to_write :  STD_LOGIC;
                signal wait_for_ext_ssram_s1_counter :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of adsc_n_to_the_ext_ssram : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of bw_n_to_the_ext_ssram : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of bwe_n_to_the_ext_ssram : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of chipenable1_n_to_the_ext_ssram : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of d1_in_a_write_cycle : signal is "FAST_OUTPUT_ENABLE_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of d1_outgoing_ext_ssram_bus_data : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of ext_ssram_bus_address : signal is "FAST_OUTPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of incoming_ext_ssram_bus_data : signal is "FAST_INPUT_REGISTER=ON";
attribute ALTERA_ATTRIBUTE of outputenable_n_to_the_ext_ssram : signal is "FAST_OUTPUT_REGISTER=ON";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT ext_ssram_bus_avalon_slave_end_xfer;
    end if;

  end process;

  ext_ssram_bus_avalon_slave_begins_xfer <= NOT d1_reasons_to_wait AND ((((internal_cpu_data_master_qualified_request_ext_ssram_s1 OR internal_cpu_instruction_master_qualified_request_ext_ssram_s1) OR internal_sgdma_rx_m_write_qualified_request_ext_ssram_s1) OR internal_sgdma_tx_m_read_qualified_request_ext_ssram_s1));
  internal_cpu_data_master_requests_ext_ssram_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(27 DOWNTO 21) & std_logic_vector'("000000000000000000000")) = std_logic_vector'("1000001000000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --~chipenable1_n_to_the_ext_ssram of type chipselect to ~p1_chipenable1_n_to_the_ext_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      chipenable1_n_to_the_ext_ssram <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      chipenable1_n_to_the_ext_ssram <= p1_chipenable1_n_to_the_ext_ssram;
    end if;

  end process;

  ext_ssram_bus_avalon_slave_write_pending <= std_logic'('0');
  --ext_ssram_bus/avalon_slave read pending calc, which is an e_assign
  ext_ssram_bus_avalon_slave_read_pending <= ((or_reduce(cpu_data_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0))) OR (or_reduce(cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0)))) OR (or_reduce(sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0)));
  --ext_ssram_bus_avalon_slave_arb_share_counter set values, which is an e_mux
  ext_ssram_bus_avalon_slave_arb_share_set_values <= std_logic'('1');
  --ext_ssram_bus_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  ext_ssram_bus_avalon_slave_non_bursting_master_requests <= ((((((((((((((internal_cpu_data_master_requests_ext_ssram_s1 OR internal_cpu_instruction_master_requests_ext_ssram_s1) OR internal_sgdma_rx_m_write_requests_ext_ssram_s1) OR internal_sgdma_tx_m_read_requests_ext_ssram_s1) OR internal_cpu_data_master_requests_ext_ssram_s1) OR internal_cpu_instruction_master_requests_ext_ssram_s1) OR internal_sgdma_rx_m_write_requests_ext_ssram_s1) OR internal_sgdma_tx_m_read_requests_ext_ssram_s1) OR internal_cpu_data_master_requests_ext_ssram_s1) OR internal_cpu_instruction_master_requests_ext_ssram_s1) OR internal_sgdma_rx_m_write_requests_ext_ssram_s1) OR internal_sgdma_tx_m_read_requests_ext_ssram_s1) OR internal_cpu_data_master_requests_ext_ssram_s1) OR internal_cpu_instruction_master_requests_ext_ssram_s1) OR internal_sgdma_rx_m_write_requests_ext_ssram_s1) OR internal_sgdma_tx_m_read_requests_ext_ssram_s1;
  --ext_ssram_bus_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  ext_ssram_bus_avalon_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --ext_ssram_bus_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  ext_ssram_bus_avalon_slave_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(ext_ssram_bus_avalon_slave_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ext_ssram_bus_avalon_slave_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(ext_ssram_bus_avalon_slave_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ext_ssram_bus_avalon_slave_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --ext_ssram_bus_avalon_slave_allgrants all slave grants, which is an e_mux
  ext_ssram_bus_avalon_slave_allgrants <= (((((((((((((((or_reduce(ext_ssram_bus_avalon_slave_grant_vector)) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector))) OR (or_reduce(ext_ssram_bus_avalon_slave_grant_vector));
  --ext_ssram_bus_avalon_slave_end_xfer assignment, which is an e_assign
  ext_ssram_bus_avalon_slave_end_xfer <= NOT ((ext_ssram_s1_waits_for_read OR ext_ssram_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave <= ext_ssram_bus_avalon_slave_end_xfer AND (((NOT ext_ssram_bus_avalon_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --ext_ssram_bus_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  ext_ssram_bus_avalon_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave AND ext_ssram_bus_avalon_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave AND NOT ext_ssram_bus_avalon_slave_non_bursting_master_requests));
  --ext_ssram_bus_avalon_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_ssram_bus_avalon_slave_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(ext_ssram_bus_avalon_slave_arb_counter_enable) = '1' then 
        ext_ssram_bus_avalon_slave_arb_share_counter <= ext_ssram_bus_avalon_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --ext_ssram_bus_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_ssram_bus_avalon_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(ext_ssram_bus_avalon_slave_master_qreq_vector) AND end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave)) OR ((end_xfer_arb_share_counter_term_ext_ssram_bus_avalon_slave AND NOT ext_ssram_bus_avalon_slave_non_bursting_master_requests)))) = '1' then 
        ext_ssram_bus_avalon_slave_slavearbiterlockenable <= ext_ssram_bus_avalon_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu/data_master ext_ssram_bus/avalon_slave arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= ext_ssram_bus_avalon_slave_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --ext_ssram_bus_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  ext_ssram_bus_avalon_slave_slavearbiterlockenable2 <= ext_ssram_bus_avalon_slave_arb_share_counter_next_value;
  --cpu/data_master ext_ssram_bus/avalon_slave arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= ext_ssram_bus_avalon_slave_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --cpu/instruction_master ext_ssram_bus/avalon_slave arbiterlock, which is an e_assign
  cpu_instruction_master_arbiterlock <= ext_ssram_bus_avalon_slave_slavearbiterlockenable AND cpu_instruction_master_continuerequest;
  --cpu/instruction_master ext_ssram_bus/avalon_slave arbiterlock2, which is an e_assign
  cpu_instruction_master_arbiterlock2 <= ext_ssram_bus_avalon_slave_slavearbiterlockenable2 AND cpu_instruction_master_continuerequest;
  --cpu/instruction_master granted ext_ssram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_instruction_master_granted_slave_ext_ssram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_instruction_master_granted_slave_ext_ssram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_instruction_master_saved_grant_ext_ssram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((ext_ssram_bus_avalon_slave_arbitration_holdoff_internal OR NOT internal_cpu_instruction_master_requests_ext_ssram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_instruction_master_granted_slave_ext_ssram_s1))))));
    end if;

  end process;

  --cpu_instruction_master_continuerequest continued request, which is an e_mux
  cpu_instruction_master_continuerequest <= (((last_cycle_cpu_instruction_master_granted_slave_ext_ssram_s1 AND internal_cpu_instruction_master_requests_ext_ssram_s1)) OR ((last_cycle_cpu_instruction_master_granted_slave_ext_ssram_s1 AND internal_cpu_instruction_master_requests_ext_ssram_s1))) OR ((last_cycle_cpu_instruction_master_granted_slave_ext_ssram_s1 AND internal_cpu_instruction_master_requests_ext_ssram_s1));
  --ext_ssram_bus_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  ext_ssram_bus_avalon_slave_any_continuerequest <= ((((((((((cpu_instruction_master_continuerequest OR sgdma_rx_m_write_continuerequest) OR sgdma_tx_m_read_continuerequest) OR cpu_data_master_continuerequest) OR sgdma_rx_m_write_continuerequest) OR sgdma_tx_m_read_continuerequest) OR cpu_data_master_continuerequest) OR cpu_instruction_master_continuerequest) OR sgdma_tx_m_read_continuerequest) OR cpu_data_master_continuerequest) OR cpu_instruction_master_continuerequest) OR sgdma_rx_m_write_continuerequest;
  --sgdma_rx/m_write ext_ssram_bus/avalon_slave arbiterlock, which is an e_assign
  sgdma_rx_m_write_arbiterlock <= ext_ssram_bus_avalon_slave_slavearbiterlockenable AND sgdma_rx_m_write_continuerequest;
  --sgdma_rx/m_write ext_ssram_bus/avalon_slave arbiterlock2, which is an e_assign
  sgdma_rx_m_write_arbiterlock2 <= ext_ssram_bus_avalon_slave_slavearbiterlockenable2 AND sgdma_rx_m_write_continuerequest;
  --sgdma_rx/m_write granted ext_ssram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_rx_m_write_granted_slave_ext_ssram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_rx_m_write_granted_slave_ext_ssram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_rx_m_write_saved_grant_ext_ssram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((ext_ssram_bus_avalon_slave_arbitration_holdoff_internal OR NOT internal_sgdma_rx_m_write_requests_ext_ssram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_rx_m_write_granted_slave_ext_ssram_s1))))));
    end if;

  end process;

  --sgdma_rx_m_write_continuerequest continued request, which is an e_mux
  sgdma_rx_m_write_continuerequest <= (((last_cycle_sgdma_rx_m_write_granted_slave_ext_ssram_s1 AND internal_sgdma_rx_m_write_requests_ext_ssram_s1)) OR ((last_cycle_sgdma_rx_m_write_granted_slave_ext_ssram_s1 AND internal_sgdma_rx_m_write_requests_ext_ssram_s1))) OR ((last_cycle_sgdma_rx_m_write_granted_slave_ext_ssram_s1 AND internal_sgdma_rx_m_write_requests_ext_ssram_s1));
  --sgdma_tx/m_read ext_ssram_bus/avalon_slave arbiterlock, which is an e_assign
  sgdma_tx_m_read_arbiterlock <= ext_ssram_bus_avalon_slave_slavearbiterlockenable AND sgdma_tx_m_read_continuerequest;
  --sgdma_tx/m_read ext_ssram_bus/avalon_slave arbiterlock2, which is an e_assign
  sgdma_tx_m_read_arbiterlock2 <= ext_ssram_bus_avalon_slave_slavearbiterlockenable2 AND sgdma_tx_m_read_continuerequest;
  --sgdma_tx/m_read granted ext_ssram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_tx_m_read_granted_slave_ext_ssram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_tx_m_read_granted_slave_ext_ssram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_tx_m_read_saved_grant_ext_ssram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((ext_ssram_bus_avalon_slave_arbitration_holdoff_internal OR NOT internal_sgdma_tx_m_read_requests_ext_ssram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_tx_m_read_granted_slave_ext_ssram_s1))))));
    end if;

  end process;

  --sgdma_tx_m_read_continuerequest continued request, which is an e_mux
  sgdma_tx_m_read_continuerequest <= (((last_cycle_sgdma_tx_m_read_granted_slave_ext_ssram_s1 AND internal_sgdma_tx_m_read_requests_ext_ssram_s1)) OR ((last_cycle_sgdma_tx_m_read_granted_slave_ext_ssram_s1 AND internal_sgdma_tx_m_read_requests_ext_ssram_s1))) OR ((last_cycle_sgdma_tx_m_read_granted_slave_ext_ssram_s1 AND internal_sgdma_tx_m_read_requests_ext_ssram_s1));
  internal_cpu_data_master_qualified_request_ext_ssram_s1 <= internal_cpu_data_master_requests_ext_ssram_s1 AND NOT (((((((cpu_data_master_read AND (((((ext_ssram_bus_avalon_slave_write_pending OR ((ext_ssram_bus_avalon_slave_read_pending AND NOT(((((or_reduce(cpu_data_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0))) OR (or_reduce(cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0)))) OR (or_reduce(sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0))))))))) OR to_std_logic(((std_logic_vector'("00000000000000000000000000000101")<(std_logic_vector'("00000000000000000000000000000") & (cpu_data_master_latency_counter)))))) OR (cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register)) OR (cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register))))) OR (((ext_ssram_bus_avalon_slave_read_pending) AND cpu_data_master_write))) OR cpu_instruction_master_arbiterlock) OR sgdma_rx_m_write_arbiterlock) OR sgdma_tx_m_read_arbiterlock));
  --cpu_data_master_read_data_valid_ext_ssram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_data_master_read_data_valid_ext_ssram_s1_shift_register_in <= (internal_cpu_data_master_granted_ext_ssram_s1 AND cpu_data_master_read) AND NOT ext_ssram_s1_waits_for_read;
  --shift register p1 cpu_data_master_read_data_valid_ext_ssram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_data_master_read_data_valid_ext_ssram_s1_shift_register <= A_EXT ((cpu_data_master_read_data_valid_ext_ssram_s1_shift_register & A_ToStdLogicVector(cpu_data_master_read_data_valid_ext_ssram_s1_shift_register_in)), 5);
  --cpu_data_master_read_data_valid_ext_ssram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_data_valid_ext_ssram_s1_shift_register <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      cpu_data_master_read_data_valid_ext_ssram_s1_shift_register <= p1_cpu_data_master_read_data_valid_ext_ssram_s1_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_data_master_read_data_valid_ext_ssram_s1, which is an e_mux
  cpu_data_master_read_data_valid_ext_ssram_s1 <= cpu_data_master_read_data_valid_ext_ssram_s1_shift_register(4);
  --ext_ssram_bus_data register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      incoming_ext_ssram_bus_data <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      incoming_ext_ssram_bus_data <= ext_ssram_bus_data;
    end if;

  end process;

  --ext_ssram_s1_with_write_latency assignment, which is an e_assign
  ext_ssram_s1_with_write_latency <= in_a_write_cycle AND ((((internal_cpu_data_master_qualified_request_ext_ssram_s1 OR internal_cpu_instruction_master_qualified_request_ext_ssram_s1) OR internal_sgdma_rx_m_write_qualified_request_ext_ssram_s1) OR internal_sgdma_tx_m_read_qualified_request_ext_ssram_s1));
  --time to write the data, which is an e_mux
  time_to_write <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((ext_ssram_s1_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'((ext_ssram_s1_with_write_latency)) = '1'), std_logic_vector'("00000000000000000000000000000001"), std_logic_vector'("00000000000000000000000000000000"))));
  --d1_outgoing_ext_ssram_bus_data register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_outgoing_ext_ssram_bus_data <= std_logic_vector'("00000000000000000000000000000000");
    elsif clk'event and clk = '1' then
      d1_outgoing_ext_ssram_bus_data <= outgoing_ext_ssram_bus_data;
    end if;

  end process;

  --write cycle delayed by 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_in_a_write_cycle <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_in_a_write_cycle <= time_to_write;
    end if;

  end process;

  --d1_outgoing_ext_ssram_bus_data tristate driver, which is an e_assign
  ext_ssram_bus_data <= A_WE_StdLogicVector((std_logic'((d1_in_a_write_cycle)) = '1'), d1_outgoing_ext_ssram_bus_data, A_REP(std_logic'('Z'), 32));
  --outgoing_ext_ssram_bus_data mux, which is an e_mux
  outgoing_ext_ssram_bus_data <= A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ext_ssram_s1)) = '1'), cpu_data_master_writedata, sgdma_rx_m_write_writedata);
  internal_cpu_instruction_master_requests_ext_ssram_s1 <= ((to_std_logic(((Std_Logic_Vector'(cpu_instruction_master_address_to_slave(27 DOWNTO 21) & std_logic_vector'("000000000000000000000")) = std_logic_vector'("1000001000000000000000000000")))) AND (cpu_instruction_master_read))) AND cpu_instruction_master_read;
  --cpu/data_master granted ext_ssram/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_data_master_granted_slave_ext_ssram_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_data_master_granted_slave_ext_ssram_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_data_master_saved_grant_ext_ssram_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((ext_ssram_bus_avalon_slave_arbitration_holdoff_internal OR NOT internal_cpu_data_master_requests_ext_ssram_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_data_master_granted_slave_ext_ssram_s1))))));
    end if;

  end process;

  --cpu_data_master_continuerequest continued request, which is an e_mux
  cpu_data_master_continuerequest <= (((last_cycle_cpu_data_master_granted_slave_ext_ssram_s1 AND internal_cpu_data_master_requests_ext_ssram_s1)) OR ((last_cycle_cpu_data_master_granted_slave_ext_ssram_s1 AND internal_cpu_data_master_requests_ext_ssram_s1))) OR ((last_cycle_cpu_data_master_granted_slave_ext_ssram_s1 AND internal_cpu_data_master_requests_ext_ssram_s1));
  internal_cpu_instruction_master_qualified_request_ext_ssram_s1 <= internal_cpu_instruction_master_requests_ext_ssram_s1 AND NOT ((((((cpu_instruction_master_read AND (((((ext_ssram_bus_avalon_slave_write_pending OR ((ext_ssram_bus_avalon_slave_read_pending AND NOT(((((or_reduce(cpu_data_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0))) OR (or_reduce(cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0)))) OR (or_reduce(sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0))))))))) OR to_std_logic(((std_logic_vector'("00000000000000000000000000000101")<(std_logic_vector'("00000000000000000000000000000") & (cpu_instruction_master_latency_counter)))))) OR (cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register)) OR (cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register))))) OR cpu_data_master_arbiterlock) OR sgdma_rx_m_write_arbiterlock) OR sgdma_tx_m_read_arbiterlock));
  --cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register_in <= (internal_cpu_instruction_master_granted_ext_ssram_s1 AND cpu_instruction_master_read) AND NOT ext_ssram_s1_waits_for_read;
  --shift register p1 cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register <= A_EXT ((cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register & A_ToStdLogicVector(cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register_in)), 5);
  --cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register <= p1_cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_instruction_master_read_data_valid_ext_ssram_s1, which is an e_mux
  cpu_instruction_master_read_data_valid_ext_ssram_s1 <= cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register(4);
  internal_sgdma_rx_m_write_requests_ext_ssram_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_rx_m_write_address_to_slave(31 DOWNTO 21) & std_logic_vector'("000000000000000000000")) = std_logic_vector'("00001000001000000000000000000000")))) AND (sgdma_rx_m_write_write))) AND sgdma_rx_m_write_write;
  internal_sgdma_rx_m_write_qualified_request_ext_ssram_s1 <= internal_sgdma_rx_m_write_requests_ext_ssram_s1 AND NOT (((((((ext_ssram_bus_avalon_slave_read_pending) AND sgdma_rx_m_write_write)) OR cpu_data_master_arbiterlock) OR cpu_instruction_master_arbiterlock) OR sgdma_tx_m_read_arbiterlock));
  internal_sgdma_tx_m_read_requests_ext_ssram_s1 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_tx_m_read_address_to_slave(31 DOWNTO 21) & std_logic_vector'("000000000000000000000")) = std_logic_vector'("00001000001000000000000000000000")))) AND (sgdma_tx_m_read_read))) AND sgdma_tx_m_read_read;
  internal_sgdma_tx_m_read_qualified_request_ext_ssram_s1 <= internal_sgdma_tx_m_read_requests_ext_ssram_s1 AND NOT ((((((sgdma_tx_m_read_read AND ((((ext_ssram_bus_avalon_slave_write_pending OR ((ext_ssram_bus_avalon_slave_read_pending AND NOT(((((or_reduce(cpu_data_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0))) OR (or_reduce(cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0)))) OR (or_reduce(sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0))))))))) OR to_std_logic(((std_logic_vector'("00000000000000000000000000000101")<(std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_m_read_latency_counter)))))) OR (sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register))))) OR cpu_data_master_arbiterlock) OR cpu_instruction_master_arbiterlock) OR sgdma_rx_m_write_arbiterlock));
  --sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register_in <= (internal_sgdma_tx_m_read_granted_ext_ssram_s1 AND sgdma_tx_m_read_read) AND NOT ext_ssram_s1_waits_for_read;
  --shift register p1 sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register <= A_EXT ((sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register & A_ToStdLogicVector(sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register_in)), 5);
  --sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register <= std_logic_vector'("00000");
    elsif clk'event and clk = '1' then
      sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register <= p1_sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register;
    end if;

  end process;

  --local readdatavalid sgdma_tx_m_read_read_data_valid_ext_ssram_s1, which is an e_mux
  sgdma_tx_m_read_read_data_valid_ext_ssram_s1 <= sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register(4);
  --allow new arb cycle for ext_ssram_bus/avalon_slave, which is an e_assign
  ext_ssram_bus_avalon_slave_allow_new_arb_cycle <= ((NOT cpu_data_master_arbiterlock AND NOT cpu_instruction_master_arbiterlock) AND NOT sgdma_rx_m_write_arbiterlock) AND NOT sgdma_tx_m_read_arbiterlock;
  --sgdma_tx/m_read assignment into master qualified-requests vector for ext_ssram/s1, which is an e_assign
  ext_ssram_bus_avalon_slave_master_qreq_vector(0) <= internal_sgdma_tx_m_read_qualified_request_ext_ssram_s1;
  --sgdma_tx/m_read grant ext_ssram/s1, which is an e_assign
  internal_sgdma_tx_m_read_granted_ext_ssram_s1 <= ext_ssram_bus_avalon_slave_grant_vector(0);
  --sgdma_tx/m_read saved-grant ext_ssram/s1, which is an e_assign
  sgdma_tx_m_read_saved_grant_ext_ssram_s1 <= ext_ssram_bus_avalon_slave_arb_winner(0) AND internal_sgdma_tx_m_read_requests_ext_ssram_s1;
  --sgdma_rx/m_write assignment into master qualified-requests vector for ext_ssram/s1, which is an e_assign
  ext_ssram_bus_avalon_slave_master_qreq_vector(1) <= internal_sgdma_rx_m_write_qualified_request_ext_ssram_s1;
  --sgdma_rx/m_write grant ext_ssram/s1, which is an e_assign
  internal_sgdma_rx_m_write_granted_ext_ssram_s1 <= ext_ssram_bus_avalon_slave_grant_vector(1);
  --sgdma_rx/m_write saved-grant ext_ssram/s1, which is an e_assign
  sgdma_rx_m_write_saved_grant_ext_ssram_s1 <= ext_ssram_bus_avalon_slave_arb_winner(1) AND internal_sgdma_rx_m_write_requests_ext_ssram_s1;
  --cpu/instruction_master assignment into master qualified-requests vector for ext_ssram/s1, which is an e_assign
  ext_ssram_bus_avalon_slave_master_qreq_vector(2) <= internal_cpu_instruction_master_qualified_request_ext_ssram_s1;
  --cpu/instruction_master grant ext_ssram/s1, which is an e_assign
  internal_cpu_instruction_master_granted_ext_ssram_s1 <= ext_ssram_bus_avalon_slave_grant_vector(2);
  --cpu/instruction_master saved-grant ext_ssram/s1, which is an e_assign
  cpu_instruction_master_saved_grant_ext_ssram_s1 <= ext_ssram_bus_avalon_slave_arb_winner(2) AND internal_cpu_instruction_master_requests_ext_ssram_s1;
  --cpu/data_master assignment into master qualified-requests vector for ext_ssram/s1, which is an e_assign
  ext_ssram_bus_avalon_slave_master_qreq_vector(3) <= internal_cpu_data_master_qualified_request_ext_ssram_s1;
  --cpu/data_master grant ext_ssram/s1, which is an e_assign
  internal_cpu_data_master_granted_ext_ssram_s1 <= ext_ssram_bus_avalon_slave_grant_vector(3);
  --cpu/data_master saved-grant ext_ssram/s1, which is an e_assign
  cpu_data_master_saved_grant_ext_ssram_s1 <= ext_ssram_bus_avalon_slave_arb_winner(3) AND internal_cpu_data_master_requests_ext_ssram_s1;
  --ext_ssram_bus/avalon_slave chosen-master double-vector, which is an e_assign
  ext_ssram_bus_avalon_slave_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((ext_ssram_bus_avalon_slave_master_qreq_vector & ext_ssram_bus_avalon_slave_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT ext_ssram_bus_avalon_slave_master_qreq_vector & NOT ext_ssram_bus_avalon_slave_master_qreq_vector))) + (std_logic_vector'("00000") & (ext_ssram_bus_avalon_slave_arb_addend))))), 8);
  --stable onehot encoding of arb winner
  ext_ssram_bus_avalon_slave_arb_winner <= A_WE_StdLogicVector((std_logic'(((ext_ssram_bus_avalon_slave_allow_new_arb_cycle AND or_reduce(ext_ssram_bus_avalon_slave_grant_vector)))) = '1'), ext_ssram_bus_avalon_slave_grant_vector, ext_ssram_bus_avalon_slave_saved_chosen_master_vector);
  --saved ext_ssram_bus_avalon_slave_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_ssram_bus_avalon_slave_saved_chosen_master_vector <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'(ext_ssram_bus_avalon_slave_allow_new_arb_cycle) = '1' then 
        ext_ssram_bus_avalon_slave_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(ext_ssram_bus_avalon_slave_grant_vector)) = '1'), ext_ssram_bus_avalon_slave_grant_vector, ext_ssram_bus_avalon_slave_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  ext_ssram_bus_avalon_slave_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((ext_ssram_bus_avalon_slave_chosen_master_double_vector(3) OR ext_ssram_bus_avalon_slave_chosen_master_double_vector(7)))) & A_ToStdLogicVector(((ext_ssram_bus_avalon_slave_chosen_master_double_vector(2) OR ext_ssram_bus_avalon_slave_chosen_master_double_vector(6)))) & A_ToStdLogicVector(((ext_ssram_bus_avalon_slave_chosen_master_double_vector(1) OR ext_ssram_bus_avalon_slave_chosen_master_double_vector(5)))) & A_ToStdLogicVector(((ext_ssram_bus_avalon_slave_chosen_master_double_vector(0) OR ext_ssram_bus_avalon_slave_chosen_master_double_vector(4)))));
  --ext_ssram_bus/avalon_slave chosen master rotated left, which is an e_assign
  ext_ssram_bus_avalon_slave_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(ext_ssram_bus_avalon_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("0000")), (std_logic_vector'("0000000000000000000000000000") & ((A_SLL(ext_ssram_bus_avalon_slave_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 4);
  --ext_ssram_bus/avalon_slave's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_ssram_bus_avalon_slave_arb_addend <= std_logic_vector'("0001");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(ext_ssram_bus_avalon_slave_grant_vector)) = '1' then 
        ext_ssram_bus_avalon_slave_arb_addend <= A_WE_StdLogicVector((std_logic'(ext_ssram_bus_avalon_slave_end_xfer) = '1'), ext_ssram_bus_avalon_slave_chosen_master_rot_left, ext_ssram_bus_avalon_slave_grant_vector);
      end if;
    end if;

  end process;

  --~adsc_n_to_the_ext_ssram of type begintransfer to ~p1_adsc_n_to_the_ext_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      adsc_n_to_the_ext_ssram <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      adsc_n_to_the_ext_ssram <= p1_adsc_n_to_the_ext_ssram;
    end if;

  end process;

  p1_adsc_n_to_the_ext_ssram <= NOT ext_ssram_bus_avalon_slave_begins_xfer;
  --~outputenable_n_to_the_ext_ssram of type outputenable to ~p1_outputenable_n_to_the_ext_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      outputenable_n_to_the_ext_ssram <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      outputenable_n_to_the_ext_ssram <= p1_outputenable_n_to_the_ext_ssram;
    end if;

  end process;

  --~p1_outputenable_n_to_the_ext_ssram assignment, which is an e_mux
  p1_outputenable_n_to_the_ext_ssram <= NOT (((((or_reduce(cpu_data_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0))) OR (or_reduce(cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0)))) OR (or_reduce(sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0)))) OR ext_ssram_s1_in_a_read_cycle));
  p1_chipenable1_n_to_the_ext_ssram <= NOT (((((((internal_cpu_data_master_granted_ext_ssram_s1 OR internal_cpu_instruction_master_granted_ext_ssram_s1) OR internal_sgdma_rx_m_write_granted_ext_ssram_s1) OR internal_sgdma_tx_m_read_granted_ext_ssram_s1) OR (or_reduce(cpu_data_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0)))) OR (or_reduce(cpu_instruction_master_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0)))) OR (or_reduce(sgdma_tx_m_read_read_data_valid_ext_ssram_s1_shift_register(2 DOWNTO 0)))));
  --ext_ssram_bus_avalon_slave_firsttransfer first transaction, which is an e_assign
  ext_ssram_bus_avalon_slave_firsttransfer <= A_WE_StdLogic((std_logic'(ext_ssram_bus_avalon_slave_begins_xfer) = '1'), ext_ssram_bus_avalon_slave_unreg_firsttransfer, ext_ssram_bus_avalon_slave_reg_firsttransfer);
  --ext_ssram_bus_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  ext_ssram_bus_avalon_slave_unreg_firsttransfer <= NOT ((ext_ssram_bus_avalon_slave_slavearbiterlockenable AND ext_ssram_bus_avalon_slave_any_continuerequest));
  --ext_ssram_bus_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_ssram_bus_avalon_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(ext_ssram_bus_avalon_slave_begins_xfer) = '1' then 
        ext_ssram_bus_avalon_slave_reg_firsttransfer <= ext_ssram_bus_avalon_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --ext_ssram_bus_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  ext_ssram_bus_avalon_slave_beginbursttransfer_internal <= ext_ssram_bus_avalon_slave_begins_xfer;
  --ext_ssram_bus_avalon_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  ext_ssram_bus_avalon_slave_arbitration_holdoff_internal <= ext_ssram_bus_avalon_slave_begins_xfer AND ext_ssram_bus_avalon_slave_firsttransfer;
  --~bwe_n_to_the_ext_ssram of type write to ~p1_bwe_n_to_the_ext_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      bwe_n_to_the_ext_ssram <= Vector_To_Std_Logic(NOT std_logic_vector'("00000000000000000000000000000000"));
    elsif clk'event and clk = '1' then
      bwe_n_to_the_ext_ssram <= p1_bwe_n_to_the_ext_ssram;
    end if;

  end process;

  --~bw_n_to_the_ext_ssram of type byteenable to ~p1_bw_n_to_the_ext_ssram, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      bw_n_to_the_ext_ssram <= A_EXT (NOT std_logic_vector'("00000000000000000000000000000000"), 4);
    elsif clk'event and clk = '1' then
      bw_n_to_the_ext_ssram <= p1_bw_n_to_the_ext_ssram;
    end if;

  end process;

  --~p1_bwe_n_to_the_ext_ssram assignment, which is an e_mux
  p1_bwe_n_to_the_ext_ssram <= NOT ((((internal_cpu_data_master_granted_ext_ssram_s1 AND cpu_data_master_write)) OR ((internal_sgdma_rx_m_write_granted_ext_ssram_s1 AND sgdma_rx_m_write_write))));
  --ext_ssram_bus_address of type address to p1_ext_ssram_bus_address, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      ext_ssram_bus_address <= std_logic_vector'("000000000000000000000");
    elsif clk'event and clk = '1' then
      ext_ssram_bus_address <= p1_ext_ssram_bus_address;
    end if;

  end process;

  --p1_ext_ssram_bus_address mux, which is an e_mux
  p1_ext_ssram_bus_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ext_ssram_s1)) = '1'), (std_logic_vector'("0000") & (cpu_data_master_address_to_slave)), A_WE_StdLogicVector((std_logic'((internal_cpu_instruction_master_granted_ext_ssram_s1)) = '1'), (std_logic_vector'("0000") & (cpu_instruction_master_address_to_slave)), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_m_write_granted_ext_ssram_s1)) = '1'), sgdma_rx_m_write_address_to_slave, sgdma_tx_m_read_address_to_slave))), 21);
  --d1_ext_ssram_bus_avalon_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_ext_ssram_bus_avalon_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_ext_ssram_bus_avalon_slave_end_xfer <= ext_ssram_bus_avalon_slave_end_xfer;
    end if;

  end process;

  --ext_ssram_s1_waits_for_read in a cycle, which is an e_mux
  ext_ssram_s1_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ext_ssram_s1_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --ext_ssram_s1_in_a_read_cycle assignment, which is an e_assign
  ext_ssram_s1_in_a_read_cycle <= (((internal_cpu_data_master_granted_ext_ssram_s1 AND cpu_data_master_read)) OR ((internal_cpu_instruction_master_granted_ext_ssram_s1 AND cpu_instruction_master_read))) OR ((internal_sgdma_tx_m_read_granted_ext_ssram_s1 AND sgdma_tx_m_read_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= ext_ssram_s1_in_a_read_cycle;
  --ext_ssram_s1_waits_for_write in a cycle, which is an e_mux
  ext_ssram_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ext_ssram_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --ext_ssram_s1_in_a_write_cycle assignment, which is an e_assign
  ext_ssram_s1_in_a_write_cycle <= ((internal_cpu_data_master_granted_ext_ssram_s1 AND cpu_data_master_write)) OR ((internal_sgdma_rx_m_write_granted_ext_ssram_s1 AND sgdma_rx_m_write_write));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= ext_ssram_s1_in_a_write_cycle;
  wait_for_ext_ssram_s1_counter <= std_logic'('0');
  --~p1_bw_n_to_the_ext_ssram byte enable port mux, which is an e_mux
  p1_bw_n_to_the_ext_ssram <= A_EXT (NOT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_ext_ssram_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_m_write_granted_ext_ssram_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (sgdma_rx_m_write_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))))), 4);
  --vhdl renameroo for output signals
  cpu_data_master_granted_ext_ssram_s1 <= internal_cpu_data_master_granted_ext_ssram_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_ext_ssram_s1 <= internal_cpu_data_master_qualified_request_ext_ssram_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_ext_ssram_s1 <= internal_cpu_data_master_requests_ext_ssram_s1;
  --vhdl renameroo for output signals
  cpu_instruction_master_granted_ext_ssram_s1 <= internal_cpu_instruction_master_granted_ext_ssram_s1;
  --vhdl renameroo for output signals
  cpu_instruction_master_qualified_request_ext_ssram_s1 <= internal_cpu_instruction_master_qualified_request_ext_ssram_s1;
  --vhdl renameroo for output signals
  cpu_instruction_master_requests_ext_ssram_s1 <= internal_cpu_instruction_master_requests_ext_ssram_s1;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_granted_ext_ssram_s1 <= internal_sgdma_rx_m_write_granted_ext_ssram_s1;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_qualified_request_ext_ssram_s1 <= internal_sgdma_rx_m_write_qualified_request_ext_ssram_s1;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_requests_ext_ssram_s1 <= internal_sgdma_rx_m_write_requests_ext_ssram_s1;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_granted_ext_ssram_s1 <= internal_sgdma_tx_m_read_granted_ext_ssram_s1;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_qualified_request_ext_ssram_s1 <= internal_sgdma_tx_m_read_qualified_request_ext_ssram_s1;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_requests_ext_ssram_s1 <= internal_sgdma_tx_m_read_requests_ext_ssram_s1;
--synthesis translate_off
    --ext_ssram/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line26 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("0000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_data_master_granted_ext_ssram_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_instruction_master_granted_ext_ssram_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(internal_sgdma_rx_m_write_granted_ext_ssram_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_m_read_granted_ext_ssram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line26, now);
          write(write_line26, string'(": "));
          write(write_line26, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line26.all);
          deallocate (write_line26);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line27 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("0000000000000000000000000000") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_data_master_saved_grant_ext_ssram_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_saved_grant_ext_ssram_s1)))))) + (std_logic_vector'("00") & (A_TOSTDLOGICVECTOR(sgdma_rx_m_write_saved_grant_ext_ssram_s1)))))) + (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(sgdma_tx_m_read_saved_grant_ext_ssram_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line27, now);
          write(write_line27, string'(": "));
          write(write_line27, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line27.all);
          deallocate (write_line27);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ext_ssram_bus_bridge_arbitrator is 
end entity ext_ssram_bus_bridge_arbitrator;


architecture europa of ext_ssram_bus_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity high_res_timer_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal high_res_timer_s1_irq : IN STD_LOGIC;
                 signal high_res_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_high_res_timer_s1_end_xfer : OUT STD_LOGIC;
                 signal high_res_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal high_res_timer_s1_chipselect : OUT STD_LOGIC;
                 signal high_res_timer_s1_irq_from_sa : OUT STD_LOGIC;
                 signal high_res_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal high_res_timer_s1_reset_n : OUT STD_LOGIC;
                 signal high_res_timer_s1_write_n : OUT STD_LOGIC;
                 signal high_res_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pipeline_bridge_m1_granted_high_res_timer_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_high_res_timer_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_high_res_timer_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_high_res_timer_s1 : OUT STD_LOGIC
              );
end entity high_res_timer_s1_arbitrator;


architecture europa of high_res_timer_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_high_res_timer_s1 :  STD_LOGIC;
                signal high_res_timer_s1_allgrants :  STD_LOGIC;
                signal high_res_timer_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal high_res_timer_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal high_res_timer_s1_any_continuerequest :  STD_LOGIC;
                signal high_res_timer_s1_arb_counter_enable :  STD_LOGIC;
                signal high_res_timer_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal high_res_timer_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal high_res_timer_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal high_res_timer_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal high_res_timer_s1_begins_xfer :  STD_LOGIC;
                signal high_res_timer_s1_end_xfer :  STD_LOGIC;
                signal high_res_timer_s1_firsttransfer :  STD_LOGIC;
                signal high_res_timer_s1_grant_vector :  STD_LOGIC;
                signal high_res_timer_s1_in_a_read_cycle :  STD_LOGIC;
                signal high_res_timer_s1_in_a_write_cycle :  STD_LOGIC;
                signal high_res_timer_s1_master_qreq_vector :  STD_LOGIC;
                signal high_res_timer_s1_non_bursting_master_requests :  STD_LOGIC;
                signal high_res_timer_s1_reg_firsttransfer :  STD_LOGIC;
                signal high_res_timer_s1_slavearbiterlockenable :  STD_LOGIC;
                signal high_res_timer_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal high_res_timer_s1_unreg_firsttransfer :  STD_LOGIC;
                signal high_res_timer_s1_waits_for_read :  STD_LOGIC;
                signal high_res_timer_s1_waits_for_write :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_high_res_timer_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_high_res_timer_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_high_res_timer_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_high_res_timer_s1 :  STD_LOGIC;
                signal shifted_address_to_high_res_timer_s1_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_high_res_timer_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT high_res_timer_s1_end_xfer;
    end if;

  end process;

  high_res_timer_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_high_res_timer_s1);
  --assign high_res_timer_s1_readdata_from_sa = high_res_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  high_res_timer_s1_readdata_from_sa <= high_res_timer_s1_readdata;
  internal_pipeline_bridge_m1_requests_high_res_timer_s1 <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1000000000001000001000000")))) AND pipeline_bridge_m1_chipselect;
  --high_res_timer_s1_arb_share_counter set values, which is an e_mux
  high_res_timer_s1_arb_share_set_values <= std_logic_vector'("001");
  --high_res_timer_s1_non_bursting_master_requests mux, which is an e_mux
  high_res_timer_s1_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_high_res_timer_s1;
  --high_res_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  high_res_timer_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --high_res_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  high_res_timer_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(high_res_timer_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (high_res_timer_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(high_res_timer_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (high_res_timer_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --high_res_timer_s1_allgrants all slave grants, which is an e_mux
  high_res_timer_s1_allgrants <= high_res_timer_s1_grant_vector;
  --high_res_timer_s1_end_xfer assignment, which is an e_assign
  high_res_timer_s1_end_xfer <= NOT ((high_res_timer_s1_waits_for_read OR high_res_timer_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_high_res_timer_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_high_res_timer_s1 <= high_res_timer_s1_end_xfer AND (((NOT high_res_timer_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --high_res_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  high_res_timer_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_high_res_timer_s1 AND high_res_timer_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_high_res_timer_s1 AND NOT high_res_timer_s1_non_bursting_master_requests));
  --high_res_timer_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      high_res_timer_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(high_res_timer_s1_arb_counter_enable) = '1' then 
        high_res_timer_s1_arb_share_counter <= high_res_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --high_res_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      high_res_timer_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((high_res_timer_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_high_res_timer_s1)) OR ((end_xfer_arb_share_counter_term_high_res_timer_s1 AND NOT high_res_timer_s1_non_bursting_master_requests)))) = '1' then 
        high_res_timer_s1_slavearbiterlockenable <= or_reduce(high_res_timer_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 high_res_timer/s1 arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= high_res_timer_s1_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --high_res_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  high_res_timer_s1_slavearbiterlockenable2 <= or_reduce(high_res_timer_s1_arb_share_counter_next_value);
  --pipeline_bridge/m1 high_res_timer/s1 arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= high_res_timer_s1_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --high_res_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  high_res_timer_s1_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_high_res_timer_s1 <= internal_pipeline_bridge_m1_requests_high_res_timer_s1 AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_high_res_timer_s1, which is an e_mux
  pipeline_bridge_m1_read_data_valid_high_res_timer_s1 <= (internal_pipeline_bridge_m1_granted_high_res_timer_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT high_res_timer_s1_waits_for_read;
  --high_res_timer_s1_writedata mux, which is an e_mux
  high_res_timer_s1_writedata <= pipeline_bridge_m1_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_high_res_timer_s1 <= internal_pipeline_bridge_m1_qualified_request_high_res_timer_s1;
  --pipeline_bridge/m1 saved-grant high_res_timer/s1, which is an e_assign
  pipeline_bridge_m1_saved_grant_high_res_timer_s1 <= internal_pipeline_bridge_m1_requests_high_res_timer_s1;
  --allow new arb cycle for high_res_timer/s1, which is an e_assign
  high_res_timer_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  high_res_timer_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  high_res_timer_s1_master_qreq_vector <= std_logic'('1');
  --high_res_timer_s1_reset_n assignment, which is an e_assign
  high_res_timer_s1_reset_n <= reset_n;
  high_res_timer_s1_chipselect <= internal_pipeline_bridge_m1_granted_high_res_timer_s1;
  --high_res_timer_s1_firsttransfer first transaction, which is an e_assign
  high_res_timer_s1_firsttransfer <= A_WE_StdLogic((std_logic'(high_res_timer_s1_begins_xfer) = '1'), high_res_timer_s1_unreg_firsttransfer, high_res_timer_s1_reg_firsttransfer);
  --high_res_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  high_res_timer_s1_unreg_firsttransfer <= NOT ((high_res_timer_s1_slavearbiterlockenable AND high_res_timer_s1_any_continuerequest));
  --high_res_timer_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      high_res_timer_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(high_res_timer_s1_begins_xfer) = '1' then 
        high_res_timer_s1_reg_firsttransfer <= high_res_timer_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --high_res_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  high_res_timer_s1_beginbursttransfer_internal <= high_res_timer_s1_begins_xfer;
  --~high_res_timer_s1_write_n assignment, which is an e_mux
  high_res_timer_s1_write_n <= NOT ((internal_pipeline_bridge_m1_granted_high_res_timer_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect))));
  shifted_address_to_high_res_timer_s1_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --high_res_timer_s1_address mux, which is an e_mux
  high_res_timer_s1_address <= A_EXT (A_SRL(shifted_address_to_high_res_timer_s1_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_high_res_timer_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_high_res_timer_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_high_res_timer_s1_end_xfer <= high_res_timer_s1_end_xfer;
    end if;

  end process;

  --high_res_timer_s1_waits_for_read in a cycle, which is an e_mux
  high_res_timer_s1_waits_for_read <= high_res_timer_s1_in_a_read_cycle AND high_res_timer_s1_begins_xfer;
  --high_res_timer_s1_in_a_read_cycle assignment, which is an e_assign
  high_res_timer_s1_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_high_res_timer_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= high_res_timer_s1_in_a_read_cycle;
  --high_res_timer_s1_waits_for_write in a cycle, which is an e_mux
  high_res_timer_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(high_res_timer_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --high_res_timer_s1_in_a_write_cycle assignment, which is an e_assign
  high_res_timer_s1_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_high_res_timer_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= high_res_timer_s1_in_a_write_cycle;
  wait_for_high_res_timer_s1_counter <= std_logic'('0');
  --assign high_res_timer_s1_irq_from_sa = high_res_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  high_res_timer_s1_irq_from_sa <= high_res_timer_s1_irq;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_high_res_timer_s1 <= internal_pipeline_bridge_m1_granted_high_res_timer_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_high_res_timer_s1 <= internal_pipeline_bridge_m1_qualified_request_high_res_timer_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_high_res_timer_s1 <= internal_pipeline_bridge_m1_requests_high_res_timer_s1;
--synthesis translate_off
    --high_res_timer/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line28 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_high_res_timer_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line28, now);
          write(write_line28, string'(": "));
          write(write_line28, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave high_res_timer/s1"));
          write(output, write_line28.all);
          deallocate (write_line28);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity interrupt_vector_interrupt_vector_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_custom_instruction_master_combo_estatus : IN STD_LOGIC;
                 signal cpu_custom_instruction_master_combo_ipending : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal interrupt_vector_interrupt_vector_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal interrupt_vector_interrupt_vector_select : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal interrupt_vector_interrupt_vector_estatus : OUT STD_LOGIC;
                 signal interrupt_vector_interrupt_vector_ipending : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal interrupt_vector_interrupt_vector_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity interrupt_vector_interrupt_vector_arbitrator;


architecture europa of interrupt_vector_interrupt_vector_arbitrator is

begin

  interrupt_vector_interrupt_vector_estatus <= cpu_custom_instruction_master_combo_estatus;
  interrupt_vector_interrupt_vector_ipending <= cpu_custom_instruction_master_combo_ipending;
  --assign interrupt_vector_interrupt_vector_result_from_sa = interrupt_vector_interrupt_vector_result so that symbol knows where to group signals which may go to master only, which is an e_assign
  interrupt_vector_interrupt_vector_result_from_sa <= interrupt_vector_interrupt_vector_result;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity jtag_uart_avalon_jtag_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                 signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC
              );
end entity jtag_uart_avalon_jtag_slave_arbitrator;


architecture europa of jtag_uart_avalon_jtag_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allgrants :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_any_continuerequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_counter_enable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_begins_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_grant_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_read_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_in_a_write_cycle :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_master_qreq_vector :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_non_bursting_master_requests :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_unreg_firsttransfer :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_read :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waits_for_write :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal shifted_address_to_jtag_uart_avalon_jtag_slave_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_jtag_uart_avalon_jtag_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  jtag_uart_avalon_jtag_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave);
  --assign jtag_uart_avalon_jtag_slave_readdata_from_sa = jtag_uart_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readdata_from_sa <= jtag_uart_avalon_jtag_slave_readdata;
  internal_pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 3) & std_logic_vector'("000")) = std_logic_vector'("1000000000001000011000000")))) AND pipeline_bridge_m1_chipselect;
  --assign jtag_uart_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_dataavailable_from_sa <= jtag_uart_avalon_jtag_slave_dataavailable;
  --assign jtag_uart_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_readyfordata_from_sa <= jtag_uart_avalon_jtag_slave_readyfordata;
  --assign jtag_uart_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= jtag_uart_avalon_jtag_slave_waitrequest;
  --jtag_uart_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  jtag_uart_avalon_jtag_slave_arb_share_set_values <= std_logic_vector'("001");
  --jtag_uart_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --jtag_uart_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(jtag_uart_avalon_jtag_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (jtag_uart_avalon_jtag_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(jtag_uart_avalon_jtag_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (jtag_uart_avalon_jtag_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --jtag_uart_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  jtag_uart_avalon_jtag_slave_allgrants <= jtag_uart_avalon_jtag_slave_grant_vector;
  --jtag_uart_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_end_xfer <= NOT ((jtag_uart_avalon_jtag_slave_waits_for_read OR jtag_uart_avalon_jtag_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave <= jtag_uart_avalon_jtag_slave_end_xfer AND (((NOT jtag_uart_avalon_jtag_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --jtag_uart_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  jtag_uart_avalon_jtag_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND jtag_uart_avalon_jtag_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests));
  --jtag_uart_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_arb_counter_enable) = '1' then 
        jtag_uart_avalon_jtag_slave_arb_share_counter <= jtag_uart_avalon_jtag_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((jtag_uart_avalon_jtag_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave)) OR ((end_xfer_arb_share_counter_term_jtag_uart_avalon_jtag_slave AND NOT jtag_uart_avalon_jtag_slave_non_bursting_master_requests)))) = '1' then 
        jtag_uart_avalon_jtag_slave_slavearbiterlockenable <= or_reduce(jtag_uart_avalon_jtag_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 jtag_uart/avalon_jtag_slave arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 <= or_reduce(jtag_uart_avalon_jtag_slave_arb_share_counter_next_value);
  --pipeline_bridge/m1 jtag_uart/avalon_jtag_slave arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= jtag_uart_avalon_jtag_slave_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --jtag_uart_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  jtag_uart_avalon_jtag_slave_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave <= internal_pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave, which is an e_mux
  pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave <= (internal_pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT jtag_uart_avalon_jtag_slave_waits_for_read;
  --jtag_uart_avalon_jtag_slave_writedata mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_writedata <= pipeline_bridge_m1_writedata;
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave <= internal_pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  --pipeline_bridge/m1 saved-grant jtag_uart/avalon_jtag_slave, which is an e_assign
  pipeline_bridge_m1_saved_grant_jtag_uart_avalon_jtag_slave <= internal_pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
  --allow new arb cycle for jtag_uart/avalon_jtag_slave, which is an e_assign
  jtag_uart_avalon_jtag_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  jtag_uart_avalon_jtag_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  jtag_uart_avalon_jtag_slave_master_qreq_vector <= std_logic'('1');
  --jtag_uart_avalon_jtag_slave_reset_n assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_reset_n <= reset_n;
  jtag_uart_avalon_jtag_slave_chipselect <= internal_pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  --jtag_uart_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_firsttransfer <= A_WE_StdLogic((std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1'), jtag_uart_avalon_jtag_slave_unreg_firsttransfer, jtag_uart_avalon_jtag_slave_reg_firsttransfer);
  --jtag_uart_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  jtag_uart_avalon_jtag_slave_unreg_firsttransfer <= NOT ((jtag_uart_avalon_jtag_slave_slavearbiterlockenable AND jtag_uart_avalon_jtag_slave_any_continuerequest));
  --jtag_uart_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      jtag_uart_avalon_jtag_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(jtag_uart_avalon_jtag_slave_begins_xfer) = '1' then 
        jtag_uart_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_avalon_jtag_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  jtag_uart_avalon_jtag_slave_beginbursttransfer_internal <= jtag_uart_avalon_jtag_slave_begins_xfer;
  --~jtag_uart_avalon_jtag_slave_read_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_read_n <= NOT ((internal_pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))));
  --~jtag_uart_avalon_jtag_slave_write_n assignment, which is an e_mux
  jtag_uart_avalon_jtag_slave_write_n <= NOT ((internal_pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect))));
  shifted_address_to_jtag_uart_avalon_jtag_slave_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --jtag_uart_avalon_jtag_slave_address mux, which is an e_mux
  jtag_uart_avalon_jtag_slave_address <= Vector_To_Std_Logic(A_SRL(shifted_address_to_jtag_uart_avalon_jtag_slave_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")));
  --d1_jtag_uart_avalon_jtag_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_jtag_uart_avalon_jtag_slave_end_xfer <= jtag_uart_avalon_jtag_slave_end_xfer;
    end if;

  end process;

  --jtag_uart_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_read <= jtag_uart_avalon_jtag_slave_in_a_read_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= jtag_uart_avalon_jtag_slave_in_a_read_cycle;
  --jtag_uart_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  jtag_uart_avalon_jtag_slave_waits_for_write <= jtag_uart_avalon_jtag_slave_in_a_write_cycle AND internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --jtag_uart_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  jtag_uart_avalon_jtag_slave_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= jtag_uart_avalon_jtag_slave_in_a_write_cycle;
  wait_for_jtag_uart_avalon_jtag_slave_counter <= std_logic'('0');
  --assign jtag_uart_avalon_jtag_slave_irq_from_sa = jtag_uart_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  jtag_uart_avalon_jtag_slave_irq_from_sa <= jtag_uart_avalon_jtag_slave_irq;
  --vhdl renameroo for output signals
  jtag_uart_avalon_jtag_slave_waitrequest_from_sa <= internal_jtag_uart_avalon_jtag_slave_waitrequest_from_sa;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave <= internal_pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave <= internal_pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave <= internal_pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave;
--synthesis translate_off
    --jtag_uart/avalon_jtag_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line29 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line29, now);
          write(write_line29, string'(": "));
          write(write_line29, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave jtag_uart/avalon_jtag_slave"));
          write(output, write_line29.all);
          deallocate (write_line29);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity lcd_display_control_slave_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal lcd_display_control_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_lcd_display_control_slave_end_xfer : OUT STD_LOGIC;
                 signal lcd_display_control_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal lcd_display_control_slave_begintransfer : OUT STD_LOGIC;
                 signal lcd_display_control_slave_read : OUT STD_LOGIC;
                 signal lcd_display_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal lcd_display_control_slave_wait_counter_eq_0 : OUT STD_LOGIC;
                 signal lcd_display_control_slave_write : OUT STD_LOGIC;
                 signal lcd_display_control_slave_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pipeline_bridge_m1_granted_lcd_display_control_slave : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_lcd_display_control_slave : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_lcd_display_control_slave : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_lcd_display_control_slave : OUT STD_LOGIC
              );
end entity lcd_display_control_slave_arbitrator;


architecture europa of lcd_display_control_slave_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_lcd_display_control_slave :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_lcd_display_control_slave_wait_counter_eq_0 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_lcd_display_control_slave :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_lcd_display_control_slave :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_lcd_display_control_slave :  STD_LOGIC;
                signal lcd_display_control_slave_allgrants :  STD_LOGIC;
                signal lcd_display_control_slave_allow_new_arb_cycle :  STD_LOGIC;
                signal lcd_display_control_slave_any_bursting_master_saved_grant :  STD_LOGIC;
                signal lcd_display_control_slave_any_continuerequest :  STD_LOGIC;
                signal lcd_display_control_slave_arb_counter_enable :  STD_LOGIC;
                signal lcd_display_control_slave_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_display_control_slave_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_display_control_slave_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal lcd_display_control_slave_beginbursttransfer_internal :  STD_LOGIC;
                signal lcd_display_control_slave_begins_xfer :  STD_LOGIC;
                signal lcd_display_control_slave_counter_load_value :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal lcd_display_control_slave_end_xfer :  STD_LOGIC;
                signal lcd_display_control_slave_firsttransfer :  STD_LOGIC;
                signal lcd_display_control_slave_grant_vector :  STD_LOGIC;
                signal lcd_display_control_slave_in_a_read_cycle :  STD_LOGIC;
                signal lcd_display_control_slave_in_a_write_cycle :  STD_LOGIC;
                signal lcd_display_control_slave_master_qreq_vector :  STD_LOGIC;
                signal lcd_display_control_slave_non_bursting_master_requests :  STD_LOGIC;
                signal lcd_display_control_slave_pretend_byte_enable :  STD_LOGIC;
                signal lcd_display_control_slave_reg_firsttransfer :  STD_LOGIC;
                signal lcd_display_control_slave_slavearbiterlockenable :  STD_LOGIC;
                signal lcd_display_control_slave_slavearbiterlockenable2 :  STD_LOGIC;
                signal lcd_display_control_slave_unreg_firsttransfer :  STD_LOGIC;
                signal lcd_display_control_slave_wait_counter :  STD_LOGIC_VECTOR (6 DOWNTO 0);
                signal lcd_display_control_slave_waits_for_read :  STD_LOGIC;
                signal lcd_display_control_slave_waits_for_write :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_lcd_display_control_slave :  STD_LOGIC;
                signal shifted_address_to_lcd_display_control_slave_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_lcd_display_control_slave_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT lcd_display_control_slave_end_xfer;
    end if;

  end process;

  lcd_display_control_slave_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_lcd_display_control_slave);
  --assign lcd_display_control_slave_readdata_from_sa = lcd_display_control_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  lcd_display_control_slave_readdata_from_sa <= lcd_display_control_slave_readdata;
  internal_pipeline_bridge_m1_requests_lcd_display_control_slave <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000000001000010000000")))) AND pipeline_bridge_m1_chipselect;
  --lcd_display_control_slave_arb_share_counter set values, which is an e_mux
  lcd_display_control_slave_arb_share_set_values <= std_logic_vector'("001");
  --lcd_display_control_slave_non_bursting_master_requests mux, which is an e_mux
  lcd_display_control_slave_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_lcd_display_control_slave;
  --lcd_display_control_slave_any_bursting_master_saved_grant mux, which is an e_mux
  lcd_display_control_slave_any_bursting_master_saved_grant <= std_logic'('0');
  --lcd_display_control_slave_arb_share_counter_next_value assignment, which is an e_assign
  lcd_display_control_slave_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(lcd_display_control_slave_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (lcd_display_control_slave_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(lcd_display_control_slave_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (lcd_display_control_slave_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --lcd_display_control_slave_allgrants all slave grants, which is an e_mux
  lcd_display_control_slave_allgrants <= lcd_display_control_slave_grant_vector;
  --lcd_display_control_slave_end_xfer assignment, which is an e_assign
  lcd_display_control_slave_end_xfer <= NOT ((lcd_display_control_slave_waits_for_read OR lcd_display_control_slave_waits_for_write));
  --end_xfer_arb_share_counter_term_lcd_display_control_slave arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_lcd_display_control_slave <= lcd_display_control_slave_end_xfer AND (((NOT lcd_display_control_slave_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --lcd_display_control_slave_arb_share_counter arbitration counter enable, which is an e_assign
  lcd_display_control_slave_arb_counter_enable <= ((end_xfer_arb_share_counter_term_lcd_display_control_slave AND lcd_display_control_slave_allgrants)) OR ((end_xfer_arb_share_counter_term_lcd_display_control_slave AND NOT lcd_display_control_slave_non_bursting_master_requests));
  --lcd_display_control_slave_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_display_control_slave_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_display_control_slave_arb_counter_enable) = '1' then 
        lcd_display_control_slave_arb_share_counter <= lcd_display_control_slave_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --lcd_display_control_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_display_control_slave_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((lcd_display_control_slave_master_qreq_vector AND end_xfer_arb_share_counter_term_lcd_display_control_slave)) OR ((end_xfer_arb_share_counter_term_lcd_display_control_slave AND NOT lcd_display_control_slave_non_bursting_master_requests)))) = '1' then 
        lcd_display_control_slave_slavearbiterlockenable <= or_reduce(lcd_display_control_slave_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 lcd_display/control_slave arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= lcd_display_control_slave_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --lcd_display_control_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  lcd_display_control_slave_slavearbiterlockenable2 <= or_reduce(lcd_display_control_slave_arb_share_counter_next_value);
  --pipeline_bridge/m1 lcd_display/control_slave arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= lcd_display_control_slave_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --lcd_display_control_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  lcd_display_control_slave_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_lcd_display_control_slave <= internal_pipeline_bridge_m1_requests_lcd_display_control_slave AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_lcd_display_control_slave, which is an e_mux
  pipeline_bridge_m1_read_data_valid_lcd_display_control_slave <= (internal_pipeline_bridge_m1_granted_lcd_display_control_slave AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT lcd_display_control_slave_waits_for_read;
  --lcd_display_control_slave_writedata mux, which is an e_mux
  lcd_display_control_slave_writedata <= pipeline_bridge_m1_writedata (7 DOWNTO 0);
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_lcd_display_control_slave <= internal_pipeline_bridge_m1_qualified_request_lcd_display_control_slave;
  --pipeline_bridge/m1 saved-grant lcd_display/control_slave, which is an e_assign
  pipeline_bridge_m1_saved_grant_lcd_display_control_slave <= internal_pipeline_bridge_m1_requests_lcd_display_control_slave;
  --allow new arb cycle for lcd_display/control_slave, which is an e_assign
  lcd_display_control_slave_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  lcd_display_control_slave_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  lcd_display_control_slave_master_qreq_vector <= std_logic'('1');
  lcd_display_control_slave_begintransfer <= lcd_display_control_slave_begins_xfer;
  --lcd_display_control_slave_firsttransfer first transaction, which is an e_assign
  lcd_display_control_slave_firsttransfer <= A_WE_StdLogic((std_logic'(lcd_display_control_slave_begins_xfer) = '1'), lcd_display_control_slave_unreg_firsttransfer, lcd_display_control_slave_reg_firsttransfer);
  --lcd_display_control_slave_unreg_firsttransfer first transaction, which is an e_assign
  lcd_display_control_slave_unreg_firsttransfer <= NOT ((lcd_display_control_slave_slavearbiterlockenable AND lcd_display_control_slave_any_continuerequest));
  --lcd_display_control_slave_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_display_control_slave_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(lcd_display_control_slave_begins_xfer) = '1' then 
        lcd_display_control_slave_reg_firsttransfer <= lcd_display_control_slave_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --lcd_display_control_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  lcd_display_control_slave_beginbursttransfer_internal <= lcd_display_control_slave_begins_xfer;
  --lcd_display_control_slave_read assignment, which is an e_mux
  lcd_display_control_slave_read <= (((internal_pipeline_bridge_m1_granted_lcd_display_control_slave AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) AND NOT lcd_display_control_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("0000000000000000000000000") & (lcd_display_control_slave_wait_counter))<std_logic_vector'("00000000000000000000000000100110"))));
  --lcd_display_control_slave_write assignment, which is an e_mux
  lcd_display_control_slave_write <= (((((internal_pipeline_bridge_m1_granted_lcd_display_control_slave AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))) AND NOT lcd_display_control_slave_begins_xfer) AND to_std_logic((((std_logic_vector'("0000000000000000000000000") & (lcd_display_control_slave_wait_counter))>=std_logic_vector'("00000000000000000000000000100110"))))) AND to_std_logic((((std_logic_vector'("0000000000000000000000000") & (lcd_display_control_slave_wait_counter))<std_logic_vector'("00000000000000000000000001001100"))))) AND lcd_display_control_slave_pretend_byte_enable;
  shifted_address_to_lcd_display_control_slave_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --lcd_display_control_slave_address mux, which is an e_mux
  lcd_display_control_slave_address <= A_EXT (A_SRL(shifted_address_to_lcd_display_control_slave_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_lcd_display_control_slave_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_lcd_display_control_slave_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_lcd_display_control_slave_end_xfer <= lcd_display_control_slave_end_xfer;
    end if;

  end process;

  --lcd_display_control_slave_waits_for_read in a cycle, which is an e_mux
  lcd_display_control_slave_waits_for_read <= lcd_display_control_slave_in_a_read_cycle AND wait_for_lcd_display_control_slave_counter;
  --lcd_display_control_slave_in_a_read_cycle assignment, which is an e_assign
  lcd_display_control_slave_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_lcd_display_control_slave AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= lcd_display_control_slave_in_a_read_cycle;
  --lcd_display_control_slave_waits_for_write in a cycle, which is an e_mux
  lcd_display_control_slave_waits_for_write <= lcd_display_control_slave_in_a_write_cycle AND wait_for_lcd_display_control_slave_counter;
  --lcd_display_control_slave_in_a_write_cycle assignment, which is an e_assign
  lcd_display_control_slave_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_lcd_display_control_slave AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= lcd_display_control_slave_in_a_write_cycle;
  internal_lcd_display_control_slave_wait_counter_eq_0 <= to_std_logic(((std_logic_vector'("0000000000000000000000000") & (lcd_display_control_slave_wait_counter)) = std_logic_vector'("00000000000000000000000000000000")));
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      lcd_display_control_slave_wait_counter <= std_logic_vector'("0000000");
    elsif clk'event and clk = '1' then
      lcd_display_control_slave_wait_counter <= lcd_display_control_slave_counter_load_value;
    end if;

  end process;

  lcd_display_control_slave_counter_load_value <= A_EXT (A_WE_StdLogicVector((std_logic'(((lcd_display_control_slave_in_a_write_cycle AND lcd_display_control_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000001110000"), A_WE_StdLogicVector((std_logic'(((lcd_display_control_slave_in_a_read_cycle AND lcd_display_control_slave_begins_xfer))) = '1'), std_logic_vector'("000000000000000000000000001001010"), A_WE_StdLogicVector((std_logic'((NOT internal_lcd_display_control_slave_wait_counter_eq_0)) = '1'), ((std_logic_vector'("00000000000000000000000000") & (lcd_display_control_slave_wait_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000")))), 7);
  wait_for_lcd_display_control_slave_counter <= lcd_display_control_slave_begins_xfer OR NOT internal_lcd_display_control_slave_wait_counter_eq_0;
  --lcd_display_control_slave_pretend_byte_enable byte enable port mux, which is an e_mux
  lcd_display_control_slave_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_m1_granted_lcd_display_control_slave)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pipeline_bridge_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  lcd_display_control_slave_wait_counter_eq_0 <= internal_lcd_display_control_slave_wait_counter_eq_0;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_lcd_display_control_slave <= internal_pipeline_bridge_m1_granted_lcd_display_control_slave;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_lcd_display_control_slave <= internal_pipeline_bridge_m1_qualified_request_lcd_display_control_slave;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_lcd_display_control_slave <= internal_pipeline_bridge_m1_requests_lcd_display_control_slave;
--synthesis translate_off
    --lcd_display/control_slave enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line30 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_lcd_display_control_slave AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line30, now);
          write(write_line30, string'(": "));
          write(write_line30, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave lcd_display/control_slave"));
          write(output, write_line30.all);
          deallocate (write_line30);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity led_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal led_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_led_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal led_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal led_pio_s1_chipselect : OUT STD_LOGIC;
                 signal led_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal led_pio_s1_reset_n : OUT STD_LOGIC;
                 signal led_pio_s1_write_n : OUT STD_LOGIC;
                 signal led_pio_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pipeline_bridge_m1_granted_led_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_led_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_led_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_led_pio_s1 : OUT STD_LOGIC
              );
end entity led_pio_s1_arbitrator;


architecture europa of led_pio_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_led_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_led_pio_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_led_pio_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_led_pio_s1 :  STD_LOGIC;
                signal led_pio_s1_allgrants :  STD_LOGIC;
                signal led_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal led_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal led_pio_s1_any_continuerequest :  STD_LOGIC;
                signal led_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal led_pio_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal led_pio_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal led_pio_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal led_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal led_pio_s1_begins_xfer :  STD_LOGIC;
                signal led_pio_s1_end_xfer :  STD_LOGIC;
                signal led_pio_s1_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_grant_vector :  STD_LOGIC;
                signal led_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal led_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal led_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal led_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal led_pio_s1_pretend_byte_enable :  STD_LOGIC;
                signal led_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal led_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal led_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal led_pio_s1_waits_for_read :  STD_LOGIC;
                signal led_pio_s1_waits_for_write :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_led_pio_s1 :  STD_LOGIC;
                signal shifted_address_to_led_pio_s1_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_led_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT led_pio_s1_end_xfer;
    end if;

  end process;

  led_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_led_pio_s1);
  --assign led_pio_s1_readdata_from_sa = led_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  led_pio_s1_readdata_from_sa <= led_pio_s1_readdata;
  internal_pipeline_bridge_m1_requests_led_pio_s1 <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000000001000010100000")))) AND pipeline_bridge_m1_chipselect;
  --led_pio_s1_arb_share_counter set values, which is an e_mux
  led_pio_s1_arb_share_set_values <= std_logic_vector'("001");
  --led_pio_s1_non_bursting_master_requests mux, which is an e_mux
  led_pio_s1_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_led_pio_s1;
  --led_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  led_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --led_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  led_pio_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(led_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (led_pio_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(led_pio_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (led_pio_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --led_pio_s1_allgrants all slave grants, which is an e_mux
  led_pio_s1_allgrants <= led_pio_s1_grant_vector;
  --led_pio_s1_end_xfer assignment, which is an e_assign
  led_pio_s1_end_xfer <= NOT ((led_pio_s1_waits_for_read OR led_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_led_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_led_pio_s1 <= led_pio_s1_end_xfer AND (((NOT led_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --led_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  led_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_led_pio_s1 AND led_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_led_pio_s1 AND NOT led_pio_s1_non_bursting_master_requests));
  --led_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(led_pio_s1_arb_counter_enable) = '1' then 
        led_pio_s1_arb_share_counter <= led_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --led_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((led_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_led_pio_s1)) OR ((end_xfer_arb_share_counter_term_led_pio_s1 AND NOT led_pio_s1_non_bursting_master_requests)))) = '1' then 
        led_pio_s1_slavearbiterlockenable <= or_reduce(led_pio_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 led_pio/s1 arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= led_pio_s1_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --led_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  led_pio_s1_slavearbiterlockenable2 <= or_reduce(led_pio_s1_arb_share_counter_next_value);
  --pipeline_bridge/m1 led_pio/s1 arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= led_pio_s1_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --led_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  led_pio_s1_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_led_pio_s1 <= internal_pipeline_bridge_m1_requests_led_pio_s1 AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_led_pio_s1, which is an e_mux
  pipeline_bridge_m1_read_data_valid_led_pio_s1 <= (internal_pipeline_bridge_m1_granted_led_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT led_pio_s1_waits_for_read;
  --led_pio_s1_writedata mux, which is an e_mux
  led_pio_s1_writedata <= pipeline_bridge_m1_writedata (7 DOWNTO 0);
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_led_pio_s1 <= internal_pipeline_bridge_m1_qualified_request_led_pio_s1;
  --pipeline_bridge/m1 saved-grant led_pio/s1, which is an e_assign
  pipeline_bridge_m1_saved_grant_led_pio_s1 <= internal_pipeline_bridge_m1_requests_led_pio_s1;
  --allow new arb cycle for led_pio/s1, which is an e_assign
  led_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  led_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  led_pio_s1_master_qreq_vector <= std_logic'('1');
  --led_pio_s1_reset_n assignment, which is an e_assign
  led_pio_s1_reset_n <= reset_n;
  led_pio_s1_chipselect <= internal_pipeline_bridge_m1_granted_led_pio_s1;
  --led_pio_s1_firsttransfer first transaction, which is an e_assign
  led_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(led_pio_s1_begins_xfer) = '1'), led_pio_s1_unreg_firsttransfer, led_pio_s1_reg_firsttransfer);
  --led_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  led_pio_s1_unreg_firsttransfer <= NOT ((led_pio_s1_slavearbiterlockenable AND led_pio_s1_any_continuerequest));
  --led_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      led_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(led_pio_s1_begins_xfer) = '1' then 
        led_pio_s1_reg_firsttransfer <= led_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --led_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  led_pio_s1_beginbursttransfer_internal <= led_pio_s1_begins_xfer;
  --~led_pio_s1_write_n assignment, which is an e_mux
  led_pio_s1_write_n <= NOT ((((internal_pipeline_bridge_m1_granted_led_pio_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))) AND led_pio_s1_pretend_byte_enable));
  shifted_address_to_led_pio_s1_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --led_pio_s1_address mux, which is an e_mux
  led_pio_s1_address <= A_EXT (A_SRL(shifted_address_to_led_pio_s1_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_led_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_led_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_led_pio_s1_end_xfer <= led_pio_s1_end_xfer;
    end if;

  end process;

  --led_pio_s1_waits_for_read in a cycle, which is an e_mux
  led_pio_s1_waits_for_read <= led_pio_s1_in_a_read_cycle AND led_pio_s1_begins_xfer;
  --led_pio_s1_in_a_read_cycle assignment, which is an e_assign
  led_pio_s1_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_led_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= led_pio_s1_in_a_read_cycle;
  --led_pio_s1_waits_for_write in a cycle, which is an e_mux
  led_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(led_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --led_pio_s1_in_a_write_cycle assignment, which is an e_assign
  led_pio_s1_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_led_pio_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= led_pio_s1_in_a_write_cycle;
  wait_for_led_pio_s1_counter <= std_logic'('0');
  --led_pio_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  led_pio_s1_pretend_byte_enable <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_pipeline_bridge_m1_granted_led_pio_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (pipeline_bridge_m1_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))));
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_led_pio_s1 <= internal_pipeline_bridge_m1_granted_led_pio_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_led_pio_s1 <= internal_pipeline_bridge_m1_qualified_request_led_pio_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_led_pio_s1 <= internal_pipeline_bridge_m1_requests_led_pio_s1;
--synthesis translate_off
    --led_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line31 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_led_pio_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line31, now);
          write(write_line31, string'(": "));
          write(write_line31, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave led_pio/s1"));
          write(output, write_line31.all);
          deallocate (write_line31);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity packet_memory_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal packet_memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_packet_memory_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_packet_memory_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_packet_memory_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_requests_packet_memory_s1 : OUT STD_LOGIC;
                 signal d1_packet_memory_s1_end_xfer : OUT STD_LOGIC;
                 signal packet_memory_s1_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal packet_memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal packet_memory_s1_chipselect : OUT STD_LOGIC;
                 signal packet_memory_s1_clken : OUT STD_LOGIC;
                 signal packet_memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal packet_memory_s1_write : OUT STD_LOGIC;
                 signal packet_memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity packet_memory_s1_arbitrator;


architecture europa of packet_memory_s1_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_packet_memory_s1_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_packet_memory_s1_shift_register_in :  STD_LOGIC;
                signal cpu_data_master_saved_grant_packet_memory_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_packet_memory_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_packet_memory_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_packet_memory_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_packet_memory_s1 :  STD_LOGIC;
                signal p1_cpu_data_master_read_data_valid_packet_memory_s1_shift_register :  STD_LOGIC;
                signal packet_memory_s1_allgrants :  STD_LOGIC;
                signal packet_memory_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal packet_memory_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal packet_memory_s1_any_continuerequest :  STD_LOGIC;
                signal packet_memory_s1_arb_counter_enable :  STD_LOGIC;
                signal packet_memory_s1_arb_share_counter :  STD_LOGIC;
                signal packet_memory_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal packet_memory_s1_arb_share_set_values :  STD_LOGIC;
                signal packet_memory_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal packet_memory_s1_begins_xfer :  STD_LOGIC;
                signal packet_memory_s1_end_xfer :  STD_LOGIC;
                signal packet_memory_s1_firsttransfer :  STD_LOGIC;
                signal packet_memory_s1_grant_vector :  STD_LOGIC;
                signal packet_memory_s1_in_a_read_cycle :  STD_LOGIC;
                signal packet_memory_s1_in_a_write_cycle :  STD_LOGIC;
                signal packet_memory_s1_master_qreq_vector :  STD_LOGIC;
                signal packet_memory_s1_non_bursting_master_requests :  STD_LOGIC;
                signal packet_memory_s1_reg_firsttransfer :  STD_LOGIC;
                signal packet_memory_s1_slavearbiterlockenable :  STD_LOGIC;
                signal packet_memory_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal packet_memory_s1_unreg_firsttransfer :  STD_LOGIC;
                signal packet_memory_s1_waits_for_read :  STD_LOGIC;
                signal packet_memory_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_packet_memory_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_packet_memory_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT packet_memory_s1_end_xfer;
    end if;

  end process;

  packet_memory_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_packet_memory_s1);
  --assign packet_memory_s1_readdata_from_sa = packet_memory_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  packet_memory_s1_readdata_from_sa <= packet_memory_s1_readdata;
  internal_cpu_data_master_requests_packet_memory_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(27 DOWNTO 16) & std_logic_vector'("0000000000000000")) = std_logic_vector'("1000010000000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --packet_memory_s1_arb_share_counter set values, which is an e_mux
  packet_memory_s1_arb_share_set_values <= std_logic'('1');
  --packet_memory_s1_non_bursting_master_requests mux, which is an e_mux
  packet_memory_s1_non_bursting_master_requests <= internal_cpu_data_master_requests_packet_memory_s1;
  --packet_memory_s1_any_bursting_master_saved_grant mux, which is an e_mux
  packet_memory_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --packet_memory_s1_arb_share_counter_next_value assignment, which is an e_assign
  packet_memory_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(packet_memory_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(packet_memory_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(packet_memory_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(packet_memory_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --packet_memory_s1_allgrants all slave grants, which is an e_mux
  packet_memory_s1_allgrants <= packet_memory_s1_grant_vector;
  --packet_memory_s1_end_xfer assignment, which is an e_assign
  packet_memory_s1_end_xfer <= NOT ((packet_memory_s1_waits_for_read OR packet_memory_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_packet_memory_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_packet_memory_s1 <= packet_memory_s1_end_xfer AND (((NOT packet_memory_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --packet_memory_s1_arb_share_counter arbitration counter enable, which is an e_assign
  packet_memory_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_packet_memory_s1 AND packet_memory_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_packet_memory_s1 AND NOT packet_memory_s1_non_bursting_master_requests));
  --packet_memory_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      packet_memory_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(packet_memory_s1_arb_counter_enable) = '1' then 
        packet_memory_s1_arb_share_counter <= packet_memory_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --packet_memory_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      packet_memory_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((packet_memory_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_packet_memory_s1)) OR ((end_xfer_arb_share_counter_term_packet_memory_s1 AND NOT packet_memory_s1_non_bursting_master_requests)))) = '1' then 
        packet_memory_s1_slavearbiterlockenable <= packet_memory_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu/data_master packet_memory/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= packet_memory_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --packet_memory_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  packet_memory_s1_slavearbiterlockenable2 <= packet_memory_s1_arb_share_counter_next_value;
  --cpu/data_master packet_memory/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= packet_memory_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --packet_memory_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  packet_memory_s1_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_packet_memory_s1 <= internal_cpu_data_master_requests_packet_memory_s1 AND NOT ((cpu_data_master_read AND (((to_std_logic(((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("00000000000000000000000000000") & (cpu_data_master_latency_counter))))) OR (cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register)) OR (cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register)))));
  --cpu_data_master_read_data_valid_packet_memory_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  cpu_data_master_read_data_valid_packet_memory_s1_shift_register_in <= (internal_cpu_data_master_granted_packet_memory_s1 AND cpu_data_master_read) AND NOT packet_memory_s1_waits_for_read;
  --shift register p1 cpu_data_master_read_data_valid_packet_memory_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_cpu_data_master_read_data_valid_packet_memory_s1_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(cpu_data_master_read_data_valid_packet_memory_s1_shift_register) & A_ToStdLogicVector(cpu_data_master_read_data_valid_packet_memory_s1_shift_register_in)));
  --cpu_data_master_read_data_valid_packet_memory_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      cpu_data_master_read_data_valid_packet_memory_s1_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      cpu_data_master_read_data_valid_packet_memory_s1_shift_register <= p1_cpu_data_master_read_data_valid_packet_memory_s1_shift_register;
    end if;

  end process;

  --local readdatavalid cpu_data_master_read_data_valid_packet_memory_s1, which is an e_mux
  cpu_data_master_read_data_valid_packet_memory_s1 <= cpu_data_master_read_data_valid_packet_memory_s1_shift_register;
  --packet_memory_s1_writedata mux, which is an e_mux
  packet_memory_s1_writedata <= cpu_data_master_writedata;
  --mux packet_memory_s1_clken, which is an e_mux
  packet_memory_s1_clken <= std_logic'('1');
  --master is always granted when requested
  internal_cpu_data_master_granted_packet_memory_s1 <= internal_cpu_data_master_qualified_request_packet_memory_s1;
  --cpu/data_master saved-grant packet_memory/s1, which is an e_assign
  cpu_data_master_saved_grant_packet_memory_s1 <= internal_cpu_data_master_requests_packet_memory_s1;
  --allow new arb cycle for packet_memory/s1, which is an e_assign
  packet_memory_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  packet_memory_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  packet_memory_s1_master_qreq_vector <= std_logic'('1');
  packet_memory_s1_chipselect <= internal_cpu_data_master_granted_packet_memory_s1;
  --packet_memory_s1_firsttransfer first transaction, which is an e_assign
  packet_memory_s1_firsttransfer <= A_WE_StdLogic((std_logic'(packet_memory_s1_begins_xfer) = '1'), packet_memory_s1_unreg_firsttransfer, packet_memory_s1_reg_firsttransfer);
  --packet_memory_s1_unreg_firsttransfer first transaction, which is an e_assign
  packet_memory_s1_unreg_firsttransfer <= NOT ((packet_memory_s1_slavearbiterlockenable AND packet_memory_s1_any_continuerequest));
  --packet_memory_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      packet_memory_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(packet_memory_s1_begins_xfer) = '1' then 
        packet_memory_s1_reg_firsttransfer <= packet_memory_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --packet_memory_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  packet_memory_s1_beginbursttransfer_internal <= packet_memory_s1_begins_xfer;
  --packet_memory_s1_write assignment, which is an e_mux
  packet_memory_s1_write <= internal_cpu_data_master_granted_packet_memory_s1 AND cpu_data_master_write;
  shifted_address_to_packet_memory_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --packet_memory_s1_address mux, which is an e_mux
  packet_memory_s1_address <= A_EXT (A_SRL(shifted_address_to_packet_memory_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 14);
  --d1_packet_memory_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_packet_memory_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_packet_memory_s1_end_xfer <= packet_memory_s1_end_xfer;
    end if;

  end process;

  --packet_memory_s1_waits_for_read in a cycle, which is an e_mux
  packet_memory_s1_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(packet_memory_s1_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --packet_memory_s1_in_a_read_cycle assignment, which is an e_assign
  packet_memory_s1_in_a_read_cycle <= internal_cpu_data_master_granted_packet_memory_s1 AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= packet_memory_s1_in_a_read_cycle;
  --packet_memory_s1_waits_for_write in a cycle, which is an e_mux
  packet_memory_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(packet_memory_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --packet_memory_s1_in_a_write_cycle assignment, which is an e_assign
  packet_memory_s1_in_a_write_cycle <= internal_cpu_data_master_granted_packet_memory_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= packet_memory_s1_in_a_write_cycle;
  wait_for_packet_memory_s1_counter <= std_logic'('0');
  --packet_memory_s1_byteenable byte enable port mux, which is an e_mux
  packet_memory_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_packet_memory_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  cpu_data_master_granted_packet_memory_s1 <= internal_cpu_data_master_granted_packet_memory_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_packet_memory_s1 <= internal_cpu_data_master_qualified_request_packet_memory_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_packet_memory_s1 <= internal_cpu_data_master_requests_packet_memory_s1;
--synthesis translate_off
    --packet_memory/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity packet_memory_s2_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal packet_memory_s2_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_m_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal sgdma_rx_m_write_write : IN STD_LOGIC;
                 signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal sgdma_tx_m_read_read : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;

              -- outputs:
                 signal d1_packet_memory_s2_end_xfer : OUT STD_LOGIC;
                 signal packet_memory_s2_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                 signal packet_memory_s2_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal packet_memory_s2_chipselect : OUT STD_LOGIC;
                 signal packet_memory_s2_clken : OUT STD_LOGIC;
                 signal packet_memory_s2_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal packet_memory_s2_write : OUT STD_LOGIC;
                 signal packet_memory_s2_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_m_write_granted_packet_memory_s2 : OUT STD_LOGIC;
                 signal sgdma_rx_m_write_qualified_request_packet_memory_s2 : OUT STD_LOGIC;
                 signal sgdma_rx_m_write_requests_packet_memory_s2 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_granted_packet_memory_s2 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_qualified_request_packet_memory_s2 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_packet_memory_s2 : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_requests_packet_memory_s2 : OUT STD_LOGIC
              );
end entity packet_memory_s2_arbitrator;


architecture europa of packet_memory_s2_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_packet_memory_s2 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_granted_packet_memory_s2 :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_qualified_request_packet_memory_s2 :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_requests_packet_memory_s2 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_granted_packet_memory_s2 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_qualified_request_packet_memory_s2 :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_requests_packet_memory_s2 :  STD_LOGIC;
                signal last_cycle_sgdma_rx_m_write_granted_slave_packet_memory_s2 :  STD_LOGIC;
                signal last_cycle_sgdma_tx_m_read_granted_slave_packet_memory_s2 :  STD_LOGIC;
                signal p1_sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register :  STD_LOGIC;
                signal packet_memory_s2_allgrants :  STD_LOGIC;
                signal packet_memory_s2_allow_new_arb_cycle :  STD_LOGIC;
                signal packet_memory_s2_any_bursting_master_saved_grant :  STD_LOGIC;
                signal packet_memory_s2_any_continuerequest :  STD_LOGIC;
                signal packet_memory_s2_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal packet_memory_s2_arb_counter_enable :  STD_LOGIC;
                signal packet_memory_s2_arb_share_counter :  STD_LOGIC;
                signal packet_memory_s2_arb_share_counter_next_value :  STD_LOGIC;
                signal packet_memory_s2_arb_share_set_values :  STD_LOGIC;
                signal packet_memory_s2_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal packet_memory_s2_arbitration_holdoff_internal :  STD_LOGIC;
                signal packet_memory_s2_beginbursttransfer_internal :  STD_LOGIC;
                signal packet_memory_s2_begins_xfer :  STD_LOGIC;
                signal packet_memory_s2_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal packet_memory_s2_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal packet_memory_s2_end_xfer :  STD_LOGIC;
                signal packet_memory_s2_firsttransfer :  STD_LOGIC;
                signal packet_memory_s2_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal packet_memory_s2_in_a_read_cycle :  STD_LOGIC;
                signal packet_memory_s2_in_a_write_cycle :  STD_LOGIC;
                signal packet_memory_s2_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal packet_memory_s2_non_bursting_master_requests :  STD_LOGIC;
                signal packet_memory_s2_reg_firsttransfer :  STD_LOGIC;
                signal packet_memory_s2_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal packet_memory_s2_slavearbiterlockenable :  STD_LOGIC;
                signal packet_memory_s2_slavearbiterlockenable2 :  STD_LOGIC;
                signal packet_memory_s2_unreg_firsttransfer :  STD_LOGIC;
                signal packet_memory_s2_waits_for_read :  STD_LOGIC;
                signal packet_memory_s2_waits_for_write :  STD_LOGIC;
                signal sgdma_rx_m_write_arbiterlock :  STD_LOGIC;
                signal sgdma_rx_m_write_arbiterlock2 :  STD_LOGIC;
                signal sgdma_rx_m_write_continuerequest :  STD_LOGIC;
                signal sgdma_rx_m_write_saved_grant_packet_memory_s2 :  STD_LOGIC;
                signal sgdma_tx_m_read_arbiterlock :  STD_LOGIC;
                signal sgdma_tx_m_read_arbiterlock2 :  STD_LOGIC;
                signal sgdma_tx_m_read_continuerequest :  STD_LOGIC;
                signal sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register :  STD_LOGIC;
                signal sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register_in :  STD_LOGIC;
                signal sgdma_tx_m_read_saved_grant_packet_memory_s2 :  STD_LOGIC;
                signal shifted_address_to_packet_memory_s2_from_sgdma_rx_m_write :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal shifted_address_to_packet_memory_s2_from_sgdma_tx_m_read :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal wait_for_packet_memory_s2_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT packet_memory_s2_end_xfer;
    end if;

  end process;

  packet_memory_s2_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_sgdma_rx_m_write_qualified_request_packet_memory_s2 OR internal_sgdma_tx_m_read_qualified_request_packet_memory_s2));
  --assign packet_memory_s2_readdata_from_sa = packet_memory_s2_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  packet_memory_s2_readdata_from_sa <= packet_memory_s2_readdata;
  internal_sgdma_rx_m_write_requests_packet_memory_s2 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_rx_m_write_address_to_slave(31 DOWNTO 16) & std_logic_vector'("0000000000000000")) = std_logic_vector'("00001000010000000000000000000000")))) AND (sgdma_rx_m_write_write))) AND sgdma_rx_m_write_write;
  --packet_memory_s2_arb_share_counter set values, which is an e_mux
  packet_memory_s2_arb_share_set_values <= std_logic'('1');
  --packet_memory_s2_non_bursting_master_requests mux, which is an e_mux
  packet_memory_s2_non_bursting_master_requests <= ((internal_sgdma_rx_m_write_requests_packet_memory_s2 OR internal_sgdma_tx_m_read_requests_packet_memory_s2) OR internal_sgdma_rx_m_write_requests_packet_memory_s2) OR internal_sgdma_tx_m_read_requests_packet_memory_s2;
  --packet_memory_s2_any_bursting_master_saved_grant mux, which is an e_mux
  packet_memory_s2_any_bursting_master_saved_grant <= std_logic'('0');
  --packet_memory_s2_arb_share_counter_next_value assignment, which is an e_assign
  packet_memory_s2_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(packet_memory_s2_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(packet_memory_s2_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(packet_memory_s2_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(packet_memory_s2_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --packet_memory_s2_allgrants all slave grants, which is an e_mux
  packet_memory_s2_allgrants <= (((or_reduce(packet_memory_s2_grant_vector)) OR (or_reduce(packet_memory_s2_grant_vector))) OR (or_reduce(packet_memory_s2_grant_vector))) OR (or_reduce(packet_memory_s2_grant_vector));
  --packet_memory_s2_end_xfer assignment, which is an e_assign
  packet_memory_s2_end_xfer <= NOT ((packet_memory_s2_waits_for_read OR packet_memory_s2_waits_for_write));
  --end_xfer_arb_share_counter_term_packet_memory_s2 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_packet_memory_s2 <= packet_memory_s2_end_xfer AND (((NOT packet_memory_s2_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --packet_memory_s2_arb_share_counter arbitration counter enable, which is an e_assign
  packet_memory_s2_arb_counter_enable <= ((end_xfer_arb_share_counter_term_packet_memory_s2 AND packet_memory_s2_allgrants)) OR ((end_xfer_arb_share_counter_term_packet_memory_s2 AND NOT packet_memory_s2_non_bursting_master_requests));
  --packet_memory_s2_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      packet_memory_s2_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(packet_memory_s2_arb_counter_enable) = '1' then 
        packet_memory_s2_arb_share_counter <= packet_memory_s2_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --packet_memory_s2_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      packet_memory_s2_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(packet_memory_s2_master_qreq_vector) AND end_xfer_arb_share_counter_term_packet_memory_s2)) OR ((end_xfer_arb_share_counter_term_packet_memory_s2 AND NOT packet_memory_s2_non_bursting_master_requests)))) = '1' then 
        packet_memory_s2_slavearbiterlockenable <= packet_memory_s2_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sgdma_rx/m_write packet_memory/s2 arbiterlock, which is an e_assign
  sgdma_rx_m_write_arbiterlock <= packet_memory_s2_slavearbiterlockenable AND sgdma_rx_m_write_continuerequest;
  --packet_memory_s2_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  packet_memory_s2_slavearbiterlockenable2 <= packet_memory_s2_arb_share_counter_next_value;
  --sgdma_rx/m_write packet_memory/s2 arbiterlock2, which is an e_assign
  sgdma_rx_m_write_arbiterlock2 <= packet_memory_s2_slavearbiterlockenable2 AND sgdma_rx_m_write_continuerequest;
  --sgdma_tx/m_read packet_memory/s2 arbiterlock, which is an e_assign
  sgdma_tx_m_read_arbiterlock <= packet_memory_s2_slavearbiterlockenable AND sgdma_tx_m_read_continuerequest;
  --sgdma_tx/m_read packet_memory/s2 arbiterlock2, which is an e_assign
  sgdma_tx_m_read_arbiterlock2 <= packet_memory_s2_slavearbiterlockenable2 AND sgdma_tx_m_read_continuerequest;
  --sgdma_tx/m_read granted packet_memory/s2 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_tx_m_read_granted_slave_packet_memory_s2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_tx_m_read_granted_slave_packet_memory_s2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_tx_m_read_saved_grant_packet_memory_s2) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((packet_memory_s2_arbitration_holdoff_internal OR NOT internal_sgdma_tx_m_read_requests_packet_memory_s2))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_tx_m_read_granted_slave_packet_memory_s2))))));
    end if;

  end process;

  --sgdma_tx_m_read_continuerequest continued request, which is an e_mux
  sgdma_tx_m_read_continuerequest <= last_cycle_sgdma_tx_m_read_granted_slave_packet_memory_s2 AND internal_sgdma_tx_m_read_requests_packet_memory_s2;
  --packet_memory_s2_any_continuerequest at least one master continues requesting, which is an e_mux
  packet_memory_s2_any_continuerequest <= sgdma_tx_m_read_continuerequest OR sgdma_rx_m_write_continuerequest;
  internal_sgdma_rx_m_write_qualified_request_packet_memory_s2 <= internal_sgdma_rx_m_write_requests_packet_memory_s2 AND NOT (sgdma_tx_m_read_arbiterlock);
  --packet_memory_s2_writedata mux, which is an e_mux
  packet_memory_s2_writedata <= sgdma_rx_m_write_writedata;
  --mux packet_memory_s2_clken, which is an e_mux
  packet_memory_s2_clken <= std_logic'('1');
  internal_sgdma_tx_m_read_requests_packet_memory_s2 <= ((to_std_logic(((Std_Logic_Vector'(sgdma_tx_m_read_address_to_slave(31 DOWNTO 16) & std_logic_vector'("0000000000000000")) = std_logic_vector'("00001000010000000000000000000000")))) AND (sgdma_tx_m_read_read))) AND sgdma_tx_m_read_read;
  --sgdma_rx/m_write granted packet_memory/s2 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_sgdma_rx_m_write_granted_slave_packet_memory_s2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_sgdma_rx_m_write_granted_slave_packet_memory_s2 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(sgdma_rx_m_write_saved_grant_packet_memory_s2) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((packet_memory_s2_arbitration_holdoff_internal OR NOT internal_sgdma_rx_m_write_requests_packet_memory_s2))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_sgdma_rx_m_write_granted_slave_packet_memory_s2))))));
    end if;

  end process;

  --sgdma_rx_m_write_continuerequest continued request, which is an e_mux
  sgdma_rx_m_write_continuerequest <= last_cycle_sgdma_rx_m_write_granted_slave_packet_memory_s2 AND internal_sgdma_rx_m_write_requests_packet_memory_s2;
  internal_sgdma_tx_m_read_qualified_request_packet_memory_s2 <= internal_sgdma_tx_m_read_requests_packet_memory_s2 AND NOT ((((sgdma_tx_m_read_read AND ((to_std_logic(((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("00000000000000000000000000000") & (sgdma_tx_m_read_latency_counter))))) OR (sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register))))) OR sgdma_rx_m_write_arbiterlock));
  --sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register_in mux for readlatency shift register, which is an e_mux
  sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register_in <= (internal_sgdma_tx_m_read_granted_packet_memory_s2 AND sgdma_tx_m_read_read) AND NOT packet_memory_s2_waits_for_read;
  --shift register p1 sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register in if flush, otherwise shift left, which is an e_mux
  p1_sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register <= Vector_To_Std_Logic(Std_Logic_Vector'(A_ToStdLogicVector(sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register) & A_ToStdLogicVector(sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register_in)));
  --sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register <= std_logic'('0');
    elsif clk'event and clk = '1' then
      sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register <= p1_sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register;
    end if;

  end process;

  --local readdatavalid sgdma_tx_m_read_read_data_valid_packet_memory_s2, which is an e_mux
  sgdma_tx_m_read_read_data_valid_packet_memory_s2 <= sgdma_tx_m_read_read_data_valid_packet_memory_s2_shift_register;
  --allow new arb cycle for packet_memory/s2, which is an e_assign
  packet_memory_s2_allow_new_arb_cycle <= NOT sgdma_rx_m_write_arbiterlock AND NOT sgdma_tx_m_read_arbiterlock;
  --sgdma_tx/m_read assignment into master qualified-requests vector for packet_memory/s2, which is an e_assign
  packet_memory_s2_master_qreq_vector(0) <= internal_sgdma_tx_m_read_qualified_request_packet_memory_s2;
  --sgdma_tx/m_read grant packet_memory/s2, which is an e_assign
  internal_sgdma_tx_m_read_granted_packet_memory_s2 <= packet_memory_s2_grant_vector(0);
  --sgdma_tx/m_read saved-grant packet_memory/s2, which is an e_assign
  sgdma_tx_m_read_saved_grant_packet_memory_s2 <= packet_memory_s2_arb_winner(0) AND internal_sgdma_tx_m_read_requests_packet_memory_s2;
  --sgdma_rx/m_write assignment into master qualified-requests vector for packet_memory/s2, which is an e_assign
  packet_memory_s2_master_qreq_vector(1) <= internal_sgdma_rx_m_write_qualified_request_packet_memory_s2;
  --sgdma_rx/m_write grant packet_memory/s2, which is an e_assign
  internal_sgdma_rx_m_write_granted_packet_memory_s2 <= packet_memory_s2_grant_vector(1);
  --sgdma_rx/m_write saved-grant packet_memory/s2, which is an e_assign
  sgdma_rx_m_write_saved_grant_packet_memory_s2 <= packet_memory_s2_arb_winner(1) AND internal_sgdma_rx_m_write_requests_packet_memory_s2;
  --packet_memory/s2 chosen-master double-vector, which is an e_assign
  packet_memory_s2_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((packet_memory_s2_master_qreq_vector & packet_memory_s2_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT packet_memory_s2_master_qreq_vector & NOT packet_memory_s2_master_qreq_vector))) + (std_logic_vector'("000") & (packet_memory_s2_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  packet_memory_s2_arb_winner <= A_WE_StdLogicVector((std_logic'(((packet_memory_s2_allow_new_arb_cycle AND or_reduce(packet_memory_s2_grant_vector)))) = '1'), packet_memory_s2_grant_vector, packet_memory_s2_saved_chosen_master_vector);
  --saved packet_memory_s2_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      packet_memory_s2_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(packet_memory_s2_allow_new_arb_cycle) = '1' then 
        packet_memory_s2_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(packet_memory_s2_grant_vector)) = '1'), packet_memory_s2_grant_vector, packet_memory_s2_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  packet_memory_s2_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((packet_memory_s2_chosen_master_double_vector(1) OR packet_memory_s2_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((packet_memory_s2_chosen_master_double_vector(0) OR packet_memory_s2_chosen_master_double_vector(2)))));
  --packet_memory/s2 chosen master rotated left, which is an e_assign
  packet_memory_s2_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(packet_memory_s2_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(packet_memory_s2_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --packet_memory/s2's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      packet_memory_s2_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(packet_memory_s2_grant_vector)) = '1' then 
        packet_memory_s2_arb_addend <= A_WE_StdLogicVector((std_logic'(packet_memory_s2_end_xfer) = '1'), packet_memory_s2_chosen_master_rot_left, packet_memory_s2_grant_vector);
      end if;
    end if;

  end process;

  packet_memory_s2_chipselect <= internal_sgdma_rx_m_write_granted_packet_memory_s2 OR internal_sgdma_tx_m_read_granted_packet_memory_s2;
  --packet_memory_s2_firsttransfer first transaction, which is an e_assign
  packet_memory_s2_firsttransfer <= A_WE_StdLogic((std_logic'(packet_memory_s2_begins_xfer) = '1'), packet_memory_s2_unreg_firsttransfer, packet_memory_s2_reg_firsttransfer);
  --packet_memory_s2_unreg_firsttransfer first transaction, which is an e_assign
  packet_memory_s2_unreg_firsttransfer <= NOT ((packet_memory_s2_slavearbiterlockenable AND packet_memory_s2_any_continuerequest));
  --packet_memory_s2_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      packet_memory_s2_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(packet_memory_s2_begins_xfer) = '1' then 
        packet_memory_s2_reg_firsttransfer <= packet_memory_s2_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --packet_memory_s2_beginbursttransfer_internal begin burst transfer, which is an e_assign
  packet_memory_s2_beginbursttransfer_internal <= packet_memory_s2_begins_xfer;
  --packet_memory_s2_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  packet_memory_s2_arbitration_holdoff_internal <= packet_memory_s2_begins_xfer AND packet_memory_s2_firsttransfer;
  --packet_memory_s2_write assignment, which is an e_mux
  packet_memory_s2_write <= internal_sgdma_rx_m_write_granted_packet_memory_s2 AND sgdma_rx_m_write_write;
  shifted_address_to_packet_memory_s2_from_sgdma_rx_m_write <= sgdma_rx_m_write_address_to_slave;
  --packet_memory_s2_address mux, which is an e_mux
  packet_memory_s2_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_m_write_granted_packet_memory_s2)) = '1'), (A_SRL(shifted_address_to_packet_memory_s2_from_sgdma_rx_m_write,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_packet_memory_s2_from_sgdma_tx_m_read,std_logic_vector'("00000000000000000000000000000010")))), 14);
  shifted_address_to_packet_memory_s2_from_sgdma_tx_m_read <= sgdma_tx_m_read_address_to_slave;
  --d1_packet_memory_s2_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_packet_memory_s2_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_packet_memory_s2_end_xfer <= packet_memory_s2_end_xfer;
    end if;

  end process;

  --packet_memory_s2_waits_for_read in a cycle, which is an e_mux
  packet_memory_s2_waits_for_read <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(packet_memory_s2_in_a_read_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --packet_memory_s2_in_a_read_cycle assignment, which is an e_assign
  packet_memory_s2_in_a_read_cycle <= internal_sgdma_tx_m_read_granted_packet_memory_s2 AND sgdma_tx_m_read_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= packet_memory_s2_in_a_read_cycle;
  --packet_memory_s2_waits_for_write in a cycle, which is an e_mux
  packet_memory_s2_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(packet_memory_s2_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --packet_memory_s2_in_a_write_cycle assignment, which is an e_assign
  packet_memory_s2_in_a_write_cycle <= internal_sgdma_rx_m_write_granted_packet_memory_s2 AND sgdma_rx_m_write_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= packet_memory_s2_in_a_write_cycle;
  wait_for_packet_memory_s2_counter <= std_logic'('0');
  --packet_memory_s2_byteenable byte enable port mux, which is an e_mux
  packet_memory_s2_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_m_write_granted_packet_memory_s2)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (sgdma_rx_m_write_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --vhdl renameroo for output signals
  sgdma_rx_m_write_granted_packet_memory_s2 <= internal_sgdma_rx_m_write_granted_packet_memory_s2;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_qualified_request_packet_memory_s2 <= internal_sgdma_rx_m_write_qualified_request_packet_memory_s2;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_requests_packet_memory_s2 <= internal_sgdma_rx_m_write_requests_packet_memory_s2;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_granted_packet_memory_s2 <= internal_sgdma_tx_m_read_granted_packet_memory_s2;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_qualified_request_packet_memory_s2 <= internal_sgdma_tx_m_read_qualified_request_packet_memory_s2;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_requests_packet_memory_s2 <= internal_sgdma_tx_m_read_requests_packet_memory_s2;
--synthesis translate_off
    --packet_memory/s2 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line32 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_sgdma_rx_m_write_granted_packet_memory_s2))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_m_read_granted_packet_memory_s2))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line32, now);
          write(write_line32, string'(": "));
          write(write_line32, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line32.all);
          deallocate (write_line32);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line33 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(sgdma_rx_m_write_saved_grant_packet_memory_s2))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(sgdma_tx_m_read_saved_grant_packet_memory_s2))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line33, now);
          write(write_line33, string'(": "));
          write(write_line33, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line33.all);
          deallocate (write_line33);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1_module;


architecture europa of rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_4;
  empty <= NOT(full_0);
  full_5 <= std_logic'('0');
  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1_module is 
        port (
              -- inputs:
                 signal clear_fifo : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal read : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sync_reset : IN STD_LOGIC;
                 signal write : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC;
                 signal empty : OUT STD_LOGIC;
                 signal fifo_contains_ones_n : OUT STD_LOGIC;
                 signal full : OUT STD_LOGIC
              );
end entity rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1_module;


architecture europa of rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1_module is
                signal full_0 :  STD_LOGIC;
                signal full_1 :  STD_LOGIC;
                signal full_2 :  STD_LOGIC;
                signal full_3 :  STD_LOGIC;
                signal full_4 :  STD_LOGIC;
                signal full_5 :  STD_LOGIC;
                signal how_many_ones :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_minus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal one_count_plus_one :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal p0_full_0 :  STD_LOGIC;
                signal p0_stage_0 :  STD_LOGIC;
                signal p1_full_1 :  STD_LOGIC;
                signal p1_stage_1 :  STD_LOGIC;
                signal p2_full_2 :  STD_LOGIC;
                signal p2_stage_2 :  STD_LOGIC;
                signal p3_full_3 :  STD_LOGIC;
                signal p3_stage_3 :  STD_LOGIC;
                signal p4_full_4 :  STD_LOGIC;
                signal p4_stage_4 :  STD_LOGIC;
                signal stage_0 :  STD_LOGIC;
                signal stage_1 :  STD_LOGIC;
                signal stage_2 :  STD_LOGIC;
                signal stage_3 :  STD_LOGIC;
                signal stage_4 :  STD_LOGIC;
                signal updated_one_count :  STD_LOGIC_VECTOR (3 DOWNTO 0);

begin

  data_out <= stage_0;
  full <= full_4;
  empty <= NOT(full_0);
  full_5 <= std_logic'('0');
  --data_4, which is an e_mux
  p4_stage_4 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_5 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, data_in);
  --data_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_4))))) = '1' then 
        if std_logic'(((sync_reset AND full_4) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_5))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_4 <= std_logic'('0');
        else
          stage_4 <= p4_stage_4;
        end if;
      end if;
    end if;

  end process;

  --control_4, which is an e_mux
  p4_full_4 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))), std_logic_vector'("00000000000000000000000000000000")));
  --control_reg_4, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_4 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_4 <= std_logic'('0');
        else
          full_4 <= p4_full_4;
        end if;
      end if;
    end if;

  end process;

  --data_3, which is an e_mux
  p3_stage_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_4 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_4);
  --data_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_3))))) = '1' then 
        if std_logic'(((sync_reset AND full_3) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_4))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_3 <= std_logic'('0');
        else
          stage_3 <= p3_stage_3;
        end if;
      end if;
    end if;

  end process;

  --control_3, which is an e_mux
  p3_full_3 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_2, full_4);
  --control_reg_3, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_3 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_3 <= std_logic'('0');
        else
          full_3 <= p3_full_3;
        end if;
      end if;
    end if;

  end process;

  --data_2, which is an e_mux
  p2_stage_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_3 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_3);
  --data_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_2))))) = '1' then 
        if std_logic'(((sync_reset AND full_2) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_3))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_2 <= std_logic'('0');
        else
          stage_2 <= p2_stage_2;
        end if;
      end if;
    end if;

  end process;

  --control_2, which is an e_mux
  p2_full_2 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_1, full_3);
  --control_reg_2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_2 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_2 <= std_logic'('0');
        else
          full_2 <= p2_full_2;
        end if;
      end if;
    end if;

  end process;

  --data_1, which is an e_mux
  p1_stage_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_2 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_2);
  --data_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_1))))) = '1' then 
        if std_logic'(((sync_reset AND full_1) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_2))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_1 <= std_logic'('0');
        else
          stage_1 <= p1_stage_1;
        end if;
      end if;
    end if;

  end process;

  --control_1, which is an e_mux
  p1_full_1 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), full_0, full_2);
  --control_reg_1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(clear_fifo) = '1' then 
          full_1 <= std_logic'('0');
        else
          full_1 <= p1_full_1;
        end if;
      end if;
    end if;

  end process;

  --data_0, which is an e_mux
  p0_stage_0 <= A_WE_StdLogic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((full_1 AND NOT clear_fifo))))) = std_logic_vector'("00000000000000000000000000000000"))), data_in, stage_1);
  --data_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      stage_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'(((sync_reset AND full_0) AND NOT((((to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1))) = std_logic_vector'("00000000000000000000000000000000")))) AND read) AND write))))) = '1' then 
          stage_0 <= std_logic'('0');
        else
          stage_0 <= p0_stage_0;
        end if;
      end if;
    end if;

  end process;

  --control_0, which is an e_mux
  p0_full_0 <= Vector_To_Std_Logic(A_WE_StdLogicVector((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((read AND NOT(write)))))) = std_logic_vector'("00000000000000000000000000000000"))), std_logic_vector'("00000000000000000000000000000001"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(full_1)))));
  --control_reg_0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      full_0 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(((clear_fifo OR ((read XOR write))) OR ((write AND NOT(full_0))))) = '1' then 
        if std_logic'((clear_fifo AND NOT write)) = '1' then 
          full_0 <= std_logic'('0');
        else
          full_0 <= p0_full_0;
        end if;
      end if;
    end if;

  end process;

  one_count_plus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) + std_logic_vector'("000000000000000000000000000000001")), 4);
  one_count_minus_one <= A_EXT (((std_logic_vector'("00000000000000000000000000000") & (how_many_ones)) - std_logic_vector'("000000000000000000000000000000001")), 4);
  --updated_one_count, which is an e_mux
  updated_one_count <= A_EXT (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND NOT(write)))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000") & (A_WE_StdLogicVector((std_logic'(((((clear_fifo OR sync_reset)) AND write))) = '1'), (std_logic_vector'("000") & (A_TOSTDLOGICVECTOR(data_in))), A_WE_StdLogicVector((std_logic'(((((read AND (data_in)) AND write) AND (stage_0)))) = '1'), how_many_ones, A_WE_StdLogicVector((std_logic'(((write AND (data_in)))) = '1'), one_count_plus_one, A_WE_StdLogicVector((std_logic'(((read AND (stage_0)))) = '1'), one_count_minus_one, how_many_ones))))))), 4);
  --counts how many ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      how_many_ones <= std_logic_vector'("0000");
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        how_many_ones <= updated_one_count;
      end if;
    end if;

  end process;

  --this fifo contains ones in the data pipeline, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      fifo_contains_ones_n <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'((((clear_fifo OR sync_reset) OR read) OR write)) = '1' then 
        fifo_contains_ones_n <= NOT (or_reduce(updated_one_count));
      end if;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pipeline_bridge_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal cpu_data_master_debugaccess : IN STD_LOGIC;
                 signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_instruction_master_read : IN STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal pipeline_bridge_s1_endofpacket : IN STD_LOGIC;
                 signal pipeline_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_s1_readdatavalid : IN STD_LOGIC;
                 signal pipeline_bridge_s1_waitrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_data_master_requests_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_granted_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_qualified_request_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register : OUT STD_LOGIC;
                 signal cpu_instruction_master_requests_pipeline_bridge_s1 : OUT STD_LOGIC;
                 signal d1_pipeline_bridge_s1_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal pipeline_bridge_s1_arbiterlock : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_arbiterlock2 : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_burstcount : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_s1_chipselect : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_debugaccess : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                 signal pipeline_bridge_s1_read : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_s1_reset_n : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_write : OUT STD_LOGIC;
                 signal pipeline_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity pipeline_bridge_s1_arbitrator;


architecture europa of pipeline_bridge_s1_arbitrator is
component rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1_module;

component rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1_module is 
           port (
                 -- inputs:
                    signal clear_fifo : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sync_reset : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC;
                    signal empty : OUT STD_LOGIC;
                    signal fifo_contains_ones_n : OUT STD_LOGIC;
                    signal full : OUT STD_LOGIC
                 );
end component rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1_module;

                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_empty_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_data_master_rdv_fifo_output_from_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_data_master_saved_grant_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock :  STD_LOGIC;
                signal cpu_instruction_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_instruction_master_continuerequest :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_instruction_master_rdv_fifo_output_from_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_instruction_master_saved_grant_pipeline_bridge_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pipeline_bridge_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_data_master_requests_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_instruction_master_granted_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_instruction_master_qualified_request_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_cpu_instruction_master_requests_pipeline_bridge_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal last_cycle_cpu_data_master_granted_slave_pipeline_bridge_s1 :  STD_LOGIC;
                signal last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_s1 :  STD_LOGIC;
                signal module_input10 :  STD_LOGIC;
                signal module_input11 :  STD_LOGIC;
                signal module_input12 :  STD_LOGIC;
                signal module_input13 :  STD_LOGIC;
                signal module_input14 :  STD_LOGIC;
                signal module_input9 :  STD_LOGIC;
                signal pipeline_bridge_s1_allgrants :  STD_LOGIC;
                signal pipeline_bridge_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pipeline_bridge_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pipeline_bridge_s1_any_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_s1_arb_addend :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_s1_arb_counter_enable :  STD_LOGIC;
                signal pipeline_bridge_s1_arb_share_counter :  STD_LOGIC;
                signal pipeline_bridge_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal pipeline_bridge_s1_arb_share_set_values :  STD_LOGIC;
                signal pipeline_bridge_s1_arb_winner :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_s1_arbitration_holdoff_internal :  STD_LOGIC;
                signal pipeline_bridge_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pipeline_bridge_s1_begins_xfer :  STD_LOGIC;
                signal pipeline_bridge_s1_chosen_master_double_vector :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pipeline_bridge_s1_chosen_master_rot_left :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_s1_end_xfer :  STD_LOGIC;
                signal pipeline_bridge_s1_firsttransfer :  STD_LOGIC;
                signal pipeline_bridge_s1_grant_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_s1_in_a_read_cycle :  STD_LOGIC;
                signal pipeline_bridge_s1_in_a_write_cycle :  STD_LOGIC;
                signal pipeline_bridge_s1_master_qreq_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_s1_move_on_to_next_transaction :  STD_LOGIC;
                signal pipeline_bridge_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pipeline_bridge_s1_readdatavalid_from_sa :  STD_LOGIC;
                signal pipeline_bridge_s1_reg_firsttransfer :  STD_LOGIC;
                signal pipeline_bridge_s1_saved_chosen_master_vector :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pipeline_bridge_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pipeline_bridge_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pipeline_bridge_s1_waits_for_read :  STD_LOGIC;
                signal pipeline_bridge_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_pipeline_bridge_s1_from_cpu_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal shifted_address_to_pipeline_bridge_s1_from_cpu_instruction_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal wait_for_pipeline_bridge_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pipeline_bridge_s1_end_xfer;
    end if;

  end process;

  pipeline_bridge_s1_begins_xfer <= NOT d1_reasons_to_wait AND ((internal_cpu_data_master_qualified_request_pipeline_bridge_s1 OR internal_cpu_instruction_master_qualified_request_pipeline_bridge_s1));
  --assign pipeline_bridge_s1_readdatavalid_from_sa = pipeline_bridge_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  pipeline_bridge_s1_readdatavalid_from_sa <= pipeline_bridge_s1_readdatavalid;
  --assign pipeline_bridge_s1_readdata_from_sa = pipeline_bridge_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pipeline_bridge_s1_readdata_from_sa <= pipeline_bridge_s1_readdata;
  internal_cpu_data_master_requests_pipeline_bridge_s1 <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(27 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("0110000000000000000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign pipeline_bridge_s1_waitrequest_from_sa = pipeline_bridge_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_pipeline_bridge_s1_waitrequest_from_sa <= pipeline_bridge_s1_waitrequest;
  --pipeline_bridge_s1_arb_share_counter set values, which is an e_mux
  pipeline_bridge_s1_arb_share_set_values <= std_logic'('1');
  --pipeline_bridge_s1_non_bursting_master_requests mux, which is an e_mux
  pipeline_bridge_s1_non_bursting_master_requests <= ((((internal_cpu_data_master_requests_pipeline_bridge_s1 OR internal_cpu_instruction_master_requests_pipeline_bridge_s1) OR internal_cpu_data_master_requests_pipeline_bridge_s1) OR internal_cpu_instruction_master_requests_pipeline_bridge_s1) OR internal_cpu_data_master_requests_pipeline_bridge_s1) OR internal_cpu_instruction_master_requests_pipeline_bridge_s1;
  --pipeline_bridge_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pipeline_bridge_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pipeline_bridge_s1_arb_share_counter_next_value assignment, which is an e_assign
  pipeline_bridge_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pipeline_bridge_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(pipeline_bridge_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --pipeline_bridge_s1_allgrants all slave grants, which is an e_mux
  pipeline_bridge_s1_allgrants <= (((((or_reduce(pipeline_bridge_s1_grant_vector)) OR (or_reduce(pipeline_bridge_s1_grant_vector))) OR (or_reduce(pipeline_bridge_s1_grant_vector))) OR (or_reduce(pipeline_bridge_s1_grant_vector))) OR (or_reduce(pipeline_bridge_s1_grant_vector))) OR (or_reduce(pipeline_bridge_s1_grant_vector));
  --pipeline_bridge_s1_end_xfer assignment, which is an e_assign
  pipeline_bridge_s1_end_xfer <= NOT ((pipeline_bridge_s1_waits_for_read OR pipeline_bridge_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pipeline_bridge_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pipeline_bridge_s1 <= pipeline_bridge_s1_end_xfer AND (((NOT pipeline_bridge_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pipeline_bridge_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pipeline_bridge_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pipeline_bridge_s1 AND pipeline_bridge_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pipeline_bridge_s1 AND NOT pipeline_bridge_s1_non_bursting_master_requests));
  --pipeline_bridge_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(pipeline_bridge_s1_arb_counter_enable) = '1' then 
        pipeline_bridge_s1_arb_share_counter <= pipeline_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pipeline_bridge_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((or_reduce(pipeline_bridge_s1_master_qreq_vector) AND end_xfer_arb_share_counter_term_pipeline_bridge_s1)) OR ((end_xfer_arb_share_counter_term_pipeline_bridge_s1 AND NOT pipeline_bridge_s1_non_bursting_master_requests)))) = '1' then 
        pipeline_bridge_s1_slavearbiterlockenable <= pipeline_bridge_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu/data_master pipeline_bridge/s1 arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= pipeline_bridge_s1_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --pipeline_bridge_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pipeline_bridge_s1_slavearbiterlockenable2 <= pipeline_bridge_s1_arb_share_counter_next_value;
  --cpu/data_master pipeline_bridge/s1 arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= pipeline_bridge_s1_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --cpu/instruction_master pipeline_bridge/s1 arbiterlock, which is an e_assign
  cpu_instruction_master_arbiterlock <= pipeline_bridge_s1_slavearbiterlockenable AND cpu_instruction_master_continuerequest;
  --cpu/instruction_master pipeline_bridge/s1 arbiterlock2, which is an e_assign
  cpu_instruction_master_arbiterlock2 <= pipeline_bridge_s1_slavearbiterlockenable2 AND cpu_instruction_master_continuerequest;
  --cpu/instruction_master granted pipeline_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_instruction_master_saved_grant_pipeline_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((pipeline_bridge_s1_arbitration_holdoff_internal OR NOT internal_cpu_instruction_master_requests_pipeline_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_s1))))));
    end if;

  end process;

  --cpu_instruction_master_continuerequest continued request, which is an e_mux
  cpu_instruction_master_continuerequest <= last_cycle_cpu_instruction_master_granted_slave_pipeline_bridge_s1 AND internal_cpu_instruction_master_requests_pipeline_bridge_s1;
  --pipeline_bridge_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  pipeline_bridge_s1_any_continuerequest <= cpu_instruction_master_continuerequest OR cpu_data_master_continuerequest;
  internal_cpu_data_master_qualified_request_pipeline_bridge_s1 <= internal_cpu_data_master_requests_pipeline_bridge_s1 AND NOT ((((cpu_data_master_read AND ((to_std_logic(((((std_logic_vector'("00000000000000000000000000000") & (cpu_data_master_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("00000000000000000000000000000") & (cpu_data_master_latency_counter)))))) OR (cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register))))) OR cpu_instruction_master_arbiterlock));
  --unique name for pipeline_bridge_s1_move_on_to_next_transaction, which is an e_assign
  pipeline_bridge_s1_move_on_to_next_transaction <= pipeline_bridge_s1_readdatavalid_from_sa;
  --rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1 : rdv_fifo_for_cpu_data_master_to_pipeline_bridge_s1_module
    port map(
      data_out => cpu_data_master_rdv_fifo_output_from_pipeline_bridge_s1,
      empty => open,
      fifo_contains_ones_n => cpu_data_master_rdv_fifo_empty_pipeline_bridge_s1,
      full => open,
      clear_fifo => module_input9,
      clk => clk,
      data_in => internal_cpu_data_master_granted_pipeline_bridge_s1,
      read => pipeline_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input10,
      write => module_input11
    );

  module_input9 <= std_logic'('0');
  module_input10 <= std_logic'('0');
  module_input11 <= in_a_read_cycle AND NOT pipeline_bridge_s1_waits_for_read;

  cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register <= NOT cpu_data_master_rdv_fifo_empty_pipeline_bridge_s1;
  --local readdatavalid cpu_data_master_read_data_valid_pipeline_bridge_s1, which is an e_mux
  cpu_data_master_read_data_valid_pipeline_bridge_s1 <= ((pipeline_bridge_s1_readdatavalid_from_sa AND cpu_data_master_rdv_fifo_output_from_pipeline_bridge_s1)) AND NOT cpu_data_master_rdv_fifo_empty_pipeline_bridge_s1;
  --pipeline_bridge_s1_writedata mux, which is an e_mux
  pipeline_bridge_s1_writedata <= cpu_data_master_writedata;
  --assign pipeline_bridge_s1_endofpacket_from_sa = pipeline_bridge_s1_endofpacket so that symbol knows where to group signals which may go to master only, which is an e_assign
  pipeline_bridge_s1_endofpacket_from_sa <= pipeline_bridge_s1_endofpacket;
  internal_cpu_instruction_master_requests_pipeline_bridge_s1 <= ((to_std_logic(((Std_Logic_Vector'(cpu_instruction_master_address_to_slave(27 DOWNTO 25) & std_logic_vector'("0000000000000000000000000")) = std_logic_vector'("0110000000000000000000000000")))) AND (cpu_instruction_master_read))) AND cpu_instruction_master_read;
  --cpu/data_master granted pipeline_bridge/s1 last time, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      last_cycle_cpu_data_master_granted_slave_pipeline_bridge_s1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      last_cycle_cpu_data_master_granted_slave_pipeline_bridge_s1 <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(cpu_data_master_saved_grant_pipeline_bridge_s1) = '1'), std_logic_vector'("00000000000000000000000000000001"), A_WE_StdLogicVector((std_logic'(((pipeline_bridge_s1_arbitration_holdoff_internal OR NOT internal_cpu_data_master_requests_pipeline_bridge_s1))) = '1'), std_logic_vector'("00000000000000000000000000000000"), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(last_cycle_cpu_data_master_granted_slave_pipeline_bridge_s1))))));
    end if;

  end process;

  --cpu_data_master_continuerequest continued request, which is an e_mux
  cpu_data_master_continuerequest <= last_cycle_cpu_data_master_granted_slave_pipeline_bridge_s1 AND internal_cpu_data_master_requests_pipeline_bridge_s1;
  internal_cpu_instruction_master_qualified_request_pipeline_bridge_s1 <= internal_cpu_instruction_master_requests_pipeline_bridge_s1 AND NOT ((((cpu_instruction_master_read AND ((to_std_logic(((((std_logic_vector'("00000000000000000000000000000") & (cpu_instruction_master_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))) OR ((std_logic_vector'("00000000000000000000000000000001")<(std_logic_vector'("00000000000000000000000000000") & (cpu_instruction_master_latency_counter)))))) OR (cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register))))) OR cpu_data_master_arbiterlock));
  --rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1 : rdv_fifo_for_cpu_instruction_master_to_pipeline_bridge_s1_module
    port map(
      data_out => cpu_instruction_master_rdv_fifo_output_from_pipeline_bridge_s1,
      empty => open,
      fifo_contains_ones_n => cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_s1,
      full => open,
      clear_fifo => module_input12,
      clk => clk,
      data_in => internal_cpu_instruction_master_granted_pipeline_bridge_s1,
      read => pipeline_bridge_s1_move_on_to_next_transaction,
      reset_n => reset_n,
      sync_reset => module_input13,
      write => module_input14
    );

  module_input12 <= std_logic'('0');
  module_input13 <= std_logic'('0');
  module_input14 <= in_a_read_cycle AND NOT pipeline_bridge_s1_waits_for_read;

  cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register <= NOT cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_s1;
  --local readdatavalid cpu_instruction_master_read_data_valid_pipeline_bridge_s1, which is an e_mux
  cpu_instruction_master_read_data_valid_pipeline_bridge_s1 <= ((pipeline_bridge_s1_readdatavalid_from_sa AND cpu_instruction_master_rdv_fifo_output_from_pipeline_bridge_s1)) AND NOT cpu_instruction_master_rdv_fifo_empty_pipeline_bridge_s1;
  --allow new arb cycle for pipeline_bridge/s1, which is an e_assign
  pipeline_bridge_s1_allow_new_arb_cycle <= NOT cpu_data_master_arbiterlock AND NOT cpu_instruction_master_arbiterlock;
  --cpu/instruction_master assignment into master qualified-requests vector for pipeline_bridge/s1, which is an e_assign
  pipeline_bridge_s1_master_qreq_vector(0) <= internal_cpu_instruction_master_qualified_request_pipeline_bridge_s1;
  --cpu/instruction_master grant pipeline_bridge/s1, which is an e_assign
  internal_cpu_instruction_master_granted_pipeline_bridge_s1 <= pipeline_bridge_s1_grant_vector(0);
  --cpu/instruction_master saved-grant pipeline_bridge/s1, which is an e_assign
  cpu_instruction_master_saved_grant_pipeline_bridge_s1 <= pipeline_bridge_s1_arb_winner(0) AND internal_cpu_instruction_master_requests_pipeline_bridge_s1;
  --cpu/data_master assignment into master qualified-requests vector for pipeline_bridge/s1, which is an e_assign
  pipeline_bridge_s1_master_qreq_vector(1) <= internal_cpu_data_master_qualified_request_pipeline_bridge_s1;
  --cpu/data_master grant pipeline_bridge/s1, which is an e_assign
  internal_cpu_data_master_granted_pipeline_bridge_s1 <= pipeline_bridge_s1_grant_vector(1);
  --cpu/data_master saved-grant pipeline_bridge/s1, which is an e_assign
  cpu_data_master_saved_grant_pipeline_bridge_s1 <= pipeline_bridge_s1_arb_winner(1) AND internal_cpu_data_master_requests_pipeline_bridge_s1;
  --pipeline_bridge/s1 chosen-master double-vector, which is an e_assign
  pipeline_bridge_s1_chosen_master_double_vector <= A_EXT (((std_logic_vector'("0") & ((pipeline_bridge_s1_master_qreq_vector & pipeline_bridge_s1_master_qreq_vector))) AND (((std_logic_vector'("0") & (Std_Logic_Vector'(NOT pipeline_bridge_s1_master_qreq_vector & NOT pipeline_bridge_s1_master_qreq_vector))) + (std_logic_vector'("000") & (pipeline_bridge_s1_arb_addend))))), 4);
  --stable onehot encoding of arb winner
  pipeline_bridge_s1_arb_winner <= A_WE_StdLogicVector((std_logic'(((pipeline_bridge_s1_allow_new_arb_cycle AND or_reduce(pipeline_bridge_s1_grant_vector)))) = '1'), pipeline_bridge_s1_grant_vector, pipeline_bridge_s1_saved_chosen_master_vector);
  --saved pipeline_bridge_s1_grant_vector, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_s1_saved_chosen_master_vector <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(pipeline_bridge_s1_allow_new_arb_cycle) = '1' then 
        pipeline_bridge_s1_saved_chosen_master_vector <= A_WE_StdLogicVector((std_logic'(or_reduce(pipeline_bridge_s1_grant_vector)) = '1'), pipeline_bridge_s1_grant_vector, pipeline_bridge_s1_saved_chosen_master_vector);
      end if;
    end if;

  end process;

  --onehot encoding of chosen master
  pipeline_bridge_s1_grant_vector <= Std_Logic_Vector'(A_ToStdLogicVector(((pipeline_bridge_s1_chosen_master_double_vector(1) OR pipeline_bridge_s1_chosen_master_double_vector(3)))) & A_ToStdLogicVector(((pipeline_bridge_s1_chosen_master_double_vector(0) OR pipeline_bridge_s1_chosen_master_double_vector(2)))));
  --pipeline_bridge/s1 chosen master rotated left, which is an e_assign
  pipeline_bridge_s1_chosen_master_rot_left <= A_EXT (A_WE_StdLogicVector((((A_SLL(pipeline_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001")))) /= std_logic_vector'("00")), (std_logic_vector'("000000000000000000000000000000") & ((A_SLL(pipeline_bridge_s1_arb_winner,std_logic_vector'("00000000000000000000000000000001"))))), std_logic_vector'("00000000000000000000000000000001")), 2);
  --pipeline_bridge/s1's addend for next-master-grant
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_s1_arb_addend <= std_logic_vector'("01");
    elsif clk'event and clk = '1' then
      if std_logic'(or_reduce(pipeline_bridge_s1_grant_vector)) = '1' then 
        pipeline_bridge_s1_arb_addend <= A_WE_StdLogicVector((std_logic'(pipeline_bridge_s1_end_xfer) = '1'), pipeline_bridge_s1_chosen_master_rot_left, pipeline_bridge_s1_grant_vector);
      end if;
    end if;

  end process;

  --pipeline_bridge_s1_reset_n assignment, which is an e_assign
  pipeline_bridge_s1_reset_n <= reset_n;
  pipeline_bridge_s1_chipselect <= internal_cpu_data_master_granted_pipeline_bridge_s1 OR internal_cpu_instruction_master_granted_pipeline_bridge_s1;
  --pipeline_bridge_s1_firsttransfer first transaction, which is an e_assign
  pipeline_bridge_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pipeline_bridge_s1_begins_xfer) = '1'), pipeline_bridge_s1_unreg_firsttransfer, pipeline_bridge_s1_reg_firsttransfer);
  --pipeline_bridge_s1_unreg_firsttransfer first transaction, which is an e_assign
  pipeline_bridge_s1_unreg_firsttransfer <= NOT ((pipeline_bridge_s1_slavearbiterlockenable AND pipeline_bridge_s1_any_continuerequest));
  --pipeline_bridge_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pipeline_bridge_s1_begins_xfer) = '1' then 
        pipeline_bridge_s1_reg_firsttransfer <= pipeline_bridge_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pipeline_bridge_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pipeline_bridge_s1_beginbursttransfer_internal <= pipeline_bridge_s1_begins_xfer;
  --pipeline_bridge_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  pipeline_bridge_s1_arbitration_holdoff_internal <= pipeline_bridge_s1_begins_xfer AND pipeline_bridge_s1_firsttransfer;
  --pipeline_bridge_s1_read assignment, which is an e_mux
  pipeline_bridge_s1_read <= ((internal_cpu_data_master_granted_pipeline_bridge_s1 AND cpu_data_master_read)) OR ((internal_cpu_instruction_master_granted_pipeline_bridge_s1 AND cpu_instruction_master_read));
  --pipeline_bridge_s1_write assignment, which is an e_mux
  pipeline_bridge_s1_write <= internal_cpu_data_master_granted_pipeline_bridge_s1 AND cpu_data_master_write;
  shifted_address_to_pipeline_bridge_s1_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --pipeline_bridge_s1_address mux, which is an e_mux
  pipeline_bridge_s1_address <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_pipeline_bridge_s1)) = '1'), (A_SRL(shifted_address_to_pipeline_bridge_s1_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(shifted_address_to_pipeline_bridge_s1_from_cpu_instruction_master,std_logic_vector'("00000000000000000000000000000010")))), 23);
  shifted_address_to_pipeline_bridge_s1_from_cpu_instruction_master <= cpu_instruction_master_address_to_slave;
  --slaveid pipeline_bridge_s1_nativeaddress nativeaddress mux, which is an e_mux
  pipeline_bridge_s1_nativeaddress <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_pipeline_bridge_s1)) = '1'), (A_SRL(cpu_data_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010"))), (A_SRL(cpu_instruction_master_address_to_slave,std_logic_vector'("00000000000000000000000000000010")))), 23);
  --d1_pipeline_bridge_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pipeline_bridge_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pipeline_bridge_s1_end_xfer <= pipeline_bridge_s1_end_xfer;
    end if;

  end process;

  --pipeline_bridge_s1_waits_for_read in a cycle, which is an e_mux
  pipeline_bridge_s1_waits_for_read <= pipeline_bridge_s1_in_a_read_cycle AND internal_pipeline_bridge_s1_waitrequest_from_sa;
  --pipeline_bridge_s1_in_a_read_cycle assignment, which is an e_assign
  pipeline_bridge_s1_in_a_read_cycle <= ((internal_cpu_data_master_granted_pipeline_bridge_s1 AND cpu_data_master_read)) OR ((internal_cpu_instruction_master_granted_pipeline_bridge_s1 AND cpu_instruction_master_read));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pipeline_bridge_s1_in_a_read_cycle;
  --pipeline_bridge_s1_waits_for_write in a cycle, which is an e_mux
  pipeline_bridge_s1_waits_for_write <= pipeline_bridge_s1_in_a_write_cycle AND internal_pipeline_bridge_s1_waitrequest_from_sa;
  --pipeline_bridge_s1_in_a_write_cycle assignment, which is an e_assign
  pipeline_bridge_s1_in_a_write_cycle <= internal_cpu_data_master_granted_pipeline_bridge_s1 AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pipeline_bridge_s1_in_a_write_cycle;
  wait_for_pipeline_bridge_s1_counter <= std_logic'('0');
  --pipeline_bridge_s1_byteenable byte enable port mux, which is an e_mux
  pipeline_bridge_s1_byteenable <= A_EXT (A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_pipeline_bridge_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000") & (cpu_data_master_byteenable)), -SIGNED(std_logic_vector'("00000000000000000000000000000001"))), 4);
  --burstcount mux, which is an e_mux
  pipeline_bridge_s1_burstcount <= std_logic'('1');
  --pipeline_bridge/s1 arbiterlock assigned from _handle_arbiterlock, which is an e_mux
  pipeline_bridge_s1_arbiterlock <= A_WE_StdLogic((std_logic'((cpu_data_master_arbiterlock)) = '1'), cpu_data_master_arbiterlock, cpu_instruction_master_arbiterlock);
  --pipeline_bridge/s1 arbiterlock2 assigned from _handle_arbiterlock2, which is an e_mux
  pipeline_bridge_s1_arbiterlock2 <= A_WE_StdLogic((std_logic'((cpu_data_master_arbiterlock2)) = '1'), cpu_data_master_arbiterlock2, cpu_instruction_master_arbiterlock2);
  --debugaccess mux, which is an e_mux
  pipeline_bridge_s1_debugaccess <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'((internal_cpu_data_master_granted_pipeline_bridge_s1)) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_data_master_debugaccess))), std_logic_vector'("00000000000000000000000000000000")));
  --vhdl renameroo for output signals
  cpu_data_master_granted_pipeline_bridge_s1 <= internal_cpu_data_master_granted_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_pipeline_bridge_s1 <= internal_cpu_data_master_qualified_request_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  cpu_data_master_requests_pipeline_bridge_s1 <= internal_cpu_data_master_requests_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  cpu_instruction_master_granted_pipeline_bridge_s1 <= internal_cpu_instruction_master_granted_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  cpu_instruction_master_qualified_request_pipeline_bridge_s1 <= internal_cpu_instruction_master_qualified_request_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  cpu_instruction_master_requests_pipeline_bridge_s1 <= internal_cpu_instruction_master_requests_pipeline_bridge_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_s1_waitrequest_from_sa <= internal_pipeline_bridge_s1_waitrequest_from_sa;
--synthesis translate_off
    --pipeline_bridge/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line34 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_data_master_granted_pipeline_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(internal_cpu_instruction_master_granted_pipeline_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line34, now);
          write(write_line34, string'(": "));
          write(write_line34, string'("> 1 of grant signals are active simultaneously"));
          write(output, write_line34.all);
          deallocate (write_line34);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --saved_grant signals are active simultaneously, which is an e_process
    process (clk)
    VARIABLE write_line35 : line;
    begin
      if clk'event and clk = '1' then
        if (std_logic_vector'("000000000000000000000000000000") & (((std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_data_master_saved_grant_pipeline_bridge_s1))) + (std_logic_vector'("0") & (A_TOSTDLOGICVECTOR(cpu_instruction_master_saved_grant_pipeline_bridge_s1))))))>std_logic_vector'("00000000000000000000000000000001") then 
          write(write_line35, now);
          write(write_line35, string'(": "));
          write(write_line35, string'("> 1 of saved_grant signals are active simultaneously"));
          write(output, write_line35.all);
          deallocate (write_line35);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity pipeline_bridge_m1_arbitrator is 
        port (
              -- inputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa : IN STD_LOGIC;
                 signal button_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer : IN STD_LOGIC;
                 signal d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer : IN STD_LOGIC;
                 signal d1_button_pio_s1_end_xfer : IN STD_LOGIC;
                 signal d1_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                 signal d1_ext_flash_enet_bus_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal d1_high_res_timer_s1_end_xfer : IN STD_LOGIC;
                 signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                 signal d1_lcd_display_control_slave_end_xfer : IN STD_LOGIC;
                 signal d1_led_pio_s1_end_xfer : IN STD_LOGIC;
                 signal d1_reconfig_request_pio_s1_end_xfer : IN STD_LOGIC;
                 signal d1_seven_seg_pio_s1_end_xfer : IN STD_LOGIC;
                 signal d1_sgdma_rx_csr_end_xfer : IN STD_LOGIC;
                 signal d1_sgdma_tx_csr_end_xfer : IN STD_LOGIC;
                 signal d1_sys_clk_timer_s1_end_xfer : IN STD_LOGIC;
                 signal d1_uart1_s1_end_xfer : IN STD_LOGIC;
                 signal ext_flash_s1_wait_counter_eq_0 : IN STD_LOGIC;
                 signal high_res_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                 signal lcd_display_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal lcd_display_control_slave_wait_counter_eq_0 : IN STD_LOGIC;
                 signal led_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pipeline_bridge_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal pipeline_bridge_m1_byteenable_ext_flash_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_button_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_ext_flash_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_high_res_timer_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_lcd_display_control_slave : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_led_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_reconfig_request_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_seven_seg_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_sgdma_rx_csr : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_sgdma_tx_csr : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_granted_uart1_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_button_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_ext_flash_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_high_res_timer_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_lcd_display_control_slave : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_led_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_sgdma_rx_csr : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_sgdma_tx_csr : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_uart1_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_button_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_ext_flash_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_high_res_timer_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_lcd_display_control_slave : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_led_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_sgdma_rx_csr : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_sgdma_tx_csr : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_uart1_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_button_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_cpu_jtag_debug_module : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_ext_flash_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_high_res_timer_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_lcd_display_control_slave : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_led_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_reconfig_request_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_seven_seg_pio_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_sgdma_rx_csr : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_sgdma_tx_csr : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_sys_clk_timer_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_requests_uart1_s1 : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reconfig_request_pio_s1_readdata_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal seven_seg_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sgdma_rx_csr_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_csr_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sys_clk_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal uart1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal pipeline_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_dbs_write_8 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal pipeline_bridge_m1_endofpacket : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal pipeline_bridge_m1_readdatavalid : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_waitrequest : OUT STD_LOGIC
              );
end entity pipeline_bridge_m1_arbitrator;


architecture europa of pipeline_bridge_m1_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal dbs_count_enable :  STD_LOGIC;
                signal dbs_counter_overflow :  STD_LOGIC;
                signal dbs_latent_8_reg_segment_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_latent_8_reg_segment_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_latent_8_reg_segment_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal dbs_rdv_count_enable :  STD_LOGIC;
                signal dbs_rdv_counter_overflow :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal internal_pipeline_bridge_m1_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_pipeline_bridge_m1_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_pipeline_bridge_m1_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal next_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal p1_dbs_latent_8_reg_segment_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_dbs_latent_8_reg_segment_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_dbs_latent_8_reg_segment_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal p1_pipeline_bridge_m1_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_m1_address_last_time :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pipeline_bridge_m1_burstcount_last_time :  STD_LOGIC;
                signal pipeline_bridge_m1_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pipeline_bridge_m1_chipselect_last_time :  STD_LOGIC;
                signal pipeline_bridge_m1_dbs_increment :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_m1_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_m1_dbs_rdv_counter_inc :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_m1_is_granted_some_slave :  STD_LOGIC;
                signal pipeline_bridge_m1_next_dbs_rdv_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_m1_read_but_no_slave_selected :  STD_LOGIC;
                signal pipeline_bridge_m1_read_last_time :  STD_LOGIC;
                signal pipeline_bridge_m1_run :  STD_LOGIC;
                signal pipeline_bridge_m1_write_last_time :  STD_LOGIC;
                signal pipeline_bridge_m1_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pre_dbs_count_enable :  STD_LOGIC;
                signal pre_flush_pipeline_bridge_m1_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal r_2 :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in OR NOT pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in OR NOT pipeline_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_chipselect)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in OR NOT pipeline_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_chipselect)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in OR NOT pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in OR NOT pipeline_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_chipselect)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in OR NOT pipeline_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_chipselect)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_button_pio_s1 OR NOT pipeline_bridge_m1_requests_button_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_button_pio_s1 OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_button_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_button_pio_s1 OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module OR NOT pipeline_bridge_m1_requests_cpu_jtag_debug_module)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_cpu_jtag_debug_module_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((((pipeline_bridge_m1_qualified_request_ext_flash_s1 OR ((((((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)) AND NOT(pipeline_bridge_m1_byteenable_ext_flash_s1)) AND internal_pipeline_bridge_m1_dbs_address(1)) AND internal_pipeline_bridge_m1_dbs_address(0)))) OR NOT pipeline_bridge_m1_requests_ext_flash_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_ext_flash_s1 OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ext_flash_s1_wait_counter_eq_0 AND NOT d1_ext_flash_enet_bus_avalon_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((internal_pipeline_bridge_m1_dbs_address(1) AND internal_pipeline_bridge_m1_dbs_address(0))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_ext_flash_s1 OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR ((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ext_flash_s1_wait_counter_eq_0 AND NOT d1_ext_flash_enet_bus_avalon_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((internal_pipeline_bridge_m1_dbs_address(1) AND internal_pipeline_bridge_m1_dbs_address(0))))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))));
  --cascaded wait assignment, which is an e_assign
  pipeline_bridge_m1_run <= (r_0 AND r_1) AND r_2;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_high_res_timer_s1 OR NOT pipeline_bridge_m1_requests_high_res_timer_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_high_res_timer_s1 OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_high_res_timer_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_high_res_timer_s1 OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave OR NOT pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave OR NOT pipeline_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_chipselect)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave OR NOT pipeline_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT jtag_uart_avalon_jtag_slave_waitrequest_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_chipselect)))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_lcd_display_control_slave OR NOT pipeline_bridge_m1_requests_lcd_display_control_slave)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_lcd_display_control_slave OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((lcd_display_control_slave_wait_counter_eq_0 AND NOT d1_lcd_display_control_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_lcd_display_control_slave OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((lcd_display_control_slave_wait_counter_eq_0 AND NOT d1_lcd_display_control_slave_end_xfer)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_led_pio_s1 OR NOT pipeline_bridge_m1_requests_led_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_led_pio_s1 OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_led_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_led_pio_s1 OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 OR NOT pipeline_bridge_m1_requests_reconfig_request_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_reconfig_request_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))));
  --r_2 master_run cascaded wait assignment, which is an e_assign
  r_2 <= Vector_To_Std_Logic((((((((((((((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 OR NOT pipeline_bridge_m1_requests_seven_seg_pio_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_seven_seg_pio_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_sgdma_rx_csr OR NOT pipeline_bridge_m1_requests_sgdma_rx_csr)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_sgdma_rx_csr OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sgdma_rx_csr_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_sgdma_rx_csr OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_sgdma_tx_csr OR NOT pipeline_bridge_m1_requests_sgdma_tx_csr)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_sgdma_tx_csr OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sgdma_tx_csr_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_sgdma_tx_csr OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 OR NOT pipeline_bridge_m1_requests_sys_clk_timer_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 OR NOT ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_sys_clk_timer_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 OR NOT ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_qualified_request_uart1_s1 OR NOT pipeline_bridge_m1_requests_uart1_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_uart1_s1 OR NOT pipeline_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_uart1_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_chipselect)))))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT pipeline_bridge_m1_qualified_request_uart1_s1 OR NOT pipeline_bridge_m1_chipselect)))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT d1_uart1_s1_end_xfer)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_chipselect)))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_pipeline_bridge_m1_address_to_slave <= pipeline_bridge_m1_address(24 DOWNTO 0);
  --pipeline_bridge_m1_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_m1_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      pipeline_bridge_m1_read_but_no_slave_selected <= (((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND pipeline_bridge_m1_run) AND NOT pipeline_bridge_m1_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  pipeline_bridge_m1_is_granted_some_slave <= (((((((((((((pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in OR pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in) OR pipeline_bridge_m1_granted_button_pio_s1) OR pipeline_bridge_m1_granted_cpu_jtag_debug_module) OR pipeline_bridge_m1_granted_ext_flash_s1) OR pipeline_bridge_m1_granted_high_res_timer_s1) OR pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave) OR pipeline_bridge_m1_granted_lcd_display_control_slave) OR pipeline_bridge_m1_granted_led_pio_s1) OR pipeline_bridge_m1_granted_reconfig_request_pio_s1) OR pipeline_bridge_m1_granted_seven_seg_pio_s1) OR pipeline_bridge_m1_granted_sgdma_rx_csr) OR pipeline_bridge_m1_granted_sgdma_tx_csr) OR pipeline_bridge_m1_granted_sys_clk_timer_s1) OR pipeline_bridge_m1_granted_uart1_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_pipeline_bridge_m1_readdatavalid <= pipeline_bridge_m1_read_data_valid_ext_flash_s1 AND dbs_rdv_counter_overflow;
  --latent slave read data valid which is not flushed, which is an e_mux
  pipeline_bridge_m1_readdatavalid <= ((((((((((((((((((((((((((((((((((((((((((pipeline_bridge_m1_read_but_no_slave_selected OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_button_pio_s1) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_high_res_timer_s1) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_lcd_display_control_slave) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_led_pio_s1) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_sgdma_rx_csr) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_sgdma_tx_csr) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1) OR pipeline_bridge_m1_read_but_no_slave_selected) OR pre_flush_pipeline_bridge_m1_readdatavalid) OR pipeline_bridge_m1_read_data_valid_uart1_s1;
  --pipeline_bridge/m1 readdata mux, which is an e_mux
  pipeline_bridge_m1_readdata <= (((((((((((((((A_REP(NOT ((pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("0000000000000000") & (NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa)))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("0000000000000000") & (NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa))))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_button_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("0000000000000000000000000000") & (button_pio_s1_readdata_from_sa))))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR cpu_jtag_debug_module_readdata_from_sa))) AND ((A_REP(NOT pipeline_bridge_m1_read_data_valid_ext_flash_s1, 32) OR Std_Logic_Vector'(incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0(7 DOWNTO 0) & dbs_latent_8_reg_segment_2 & dbs_latent_8_reg_segment_1 & dbs_latent_8_reg_segment_0)))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_high_res_timer_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("0000000000000000") & (high_res_timer_s1_readdata_from_sa))))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR jtag_uart_avalon_jtag_slave_readdata_from_sa))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_lcd_display_control_slave AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("000000000000000000000000") & (lcd_display_control_slave_readdata_from_sa))))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_led_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("000000000000000000000000") & (led_pio_s1_readdata_from_sa))))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(reconfig_request_pio_s1_readdata_from_sa)))))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("0000000000000000") & (seven_seg_pio_s1_readdata_from_sa))))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_sgdma_rx_csr AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR sgdma_rx_csr_readdata_from_sa))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_sgdma_tx_csr AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR sgdma_tx_csr_readdata_from_sa))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("0000000000000000") & (sys_clk_timer_s1_readdata_from_sa))))) AND ((A_REP(NOT ((pipeline_bridge_m1_qualified_request_uart1_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))) , 32) OR (std_logic_vector'("0000000000000000") & (uart1_s1_readdata_from_sa))));
  --actual waitrequest port, which is an e_assign
  internal_pipeline_bridge_m1_waitrequest <= NOT pipeline_bridge_m1_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pipeline_bridge_m1_latency_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      internal_pipeline_bridge_m1_latency_counter <= p1_pipeline_bridge_m1_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_pipeline_bridge_m1_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((pipeline_bridge_m1_run AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))))) = '1'), (std_logic_vector'("0000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00")), ((std_logic_vector'("0000000000000000000000000000000") & (internal_pipeline_bridge_m1_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 2);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT (((std_logic_vector'("000000000000000000000000000000") & (A_REP(pipeline_bridge_m1_requests_ext_flash_s1, 2))) AND std_logic_vector'("00000000000000000000000000000010")), 2);
  --mux pipeline_bridge_m1_endofpacket, which is an e_mux
  pipeline_bridge_m1_endofpacket <= A_WE_StdLogic((std_logic'((pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in)) = '1'), NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa, NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa);
  --pre dbs count enable, which is an e_mux
  pre_dbs_count_enable <= Vector_To_Std_Logic((((((((NOT std_logic_vector'("00000000000000000000000000000000")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_requests_ext_flash_s1)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT(pipeline_bridge_m1_byteenable_ext_flash_s1)))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pipeline_bridge_m1_granted_ext_flash_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)))))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ext_flash_s1_wait_counter_eq_0 AND NOT d1_ext_flash_enet_bus_avalon_slave_end_xfer)))))))) OR (((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((pipeline_bridge_m1_granted_ext_flash_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))))) AND std_logic_vector'("00000000000000000000000000000001")) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((ext_flash_s1_wait_counter_eq_0 AND NOT d1_ext_flash_enet_bus_avalon_slave_end_xfer)))))))));
  --input to latent dbs-8 stored 0, which is an e_mux
  p1_dbs_latent_8_reg_segment_0 <= incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0;
  --dbs register for latent dbs-8 segment 0, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_8_reg_segment_0 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((pipeline_bridge_m1_dbs_rdv_counter(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000000")))))) = '1' then 
        dbs_latent_8_reg_segment_0 <= p1_dbs_latent_8_reg_segment_0;
      end if;
    end if;

  end process;

  --input to latent dbs-8 stored 1, which is an e_mux
  p1_dbs_latent_8_reg_segment_1 <= incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0;
  --dbs register for latent dbs-8 segment 1, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_8_reg_segment_1 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((pipeline_bridge_m1_dbs_rdv_counter(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000001")))))) = '1' then 
        dbs_latent_8_reg_segment_1 <= p1_dbs_latent_8_reg_segment_1;
      end if;
    end if;

  end process;

  --input to latent dbs-8 stored 2, which is an e_mux
  p1_dbs_latent_8_reg_segment_2 <= incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0;
  --dbs register for latent dbs-8 segment 2, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      dbs_latent_8_reg_segment_2 <= std_logic_vector'("00000000");
    elsif clk'event and clk = '1' then
      if std_logic'((dbs_rdv_count_enable AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & ((pipeline_bridge_m1_dbs_rdv_counter(1 DOWNTO 0)))) = std_logic_vector'("00000000000000000000000000000010")))))) = '1' then 
        dbs_latent_8_reg_segment_2 <= p1_dbs_latent_8_reg_segment_2;
      end if;
    end if;

  end process;

  --mux write dbs 2, which is an e_mux
  pipeline_bridge_m1_dbs_write_8 <= A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_pipeline_bridge_m1_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000000"))), pipeline_bridge_m1_writedata(7 DOWNTO 0), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_pipeline_bridge_m1_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000001"))), pipeline_bridge_m1_writedata(15 DOWNTO 8), A_WE_StdLogicVector((((std_logic_vector'("000000000000000000000000000000") & (internal_pipeline_bridge_m1_dbs_address(1 DOWNTO 0))) = std_logic_vector'("00000000000000000000000000000010"))), pipeline_bridge_m1_writedata(23 DOWNTO 16), pipeline_bridge_m1_writedata(31 DOWNTO 24))));
  --dbs count increment, which is an e_mux
  pipeline_bridge_m1_dbs_increment <= A_EXT (A_WE_StdLogicVector((std_logic'((pipeline_bridge_m1_requests_ext_flash_s1)) = '1'), std_logic_vector'("00000000000000000000000000000001"), std_logic_vector'("00000000000000000000000000000000")), 2);
  --dbs counter overflow, which is an e_assign
  dbs_counter_overflow <= internal_pipeline_bridge_m1_dbs_address(1) AND NOT((next_dbs_address(1)));
  --next master address, which is an e_assign
  next_dbs_address <= A_EXT (((std_logic_vector'("0") & (internal_pipeline_bridge_m1_dbs_address)) + (std_logic_vector'("0") & (pipeline_bridge_m1_dbs_increment))), 2);
  --dbs count enable, which is an e_mux
  dbs_count_enable <= pre_dbs_count_enable;
  --dbs counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_pipeline_bridge_m1_dbs_address <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_count_enable) = '1' then 
        internal_pipeline_bridge_m1_dbs_address <= next_dbs_address;
      end if;
    end if;

  end process;

  --p1 dbs rdv counter, which is an e_assign
  pipeline_bridge_m1_next_dbs_rdv_counter <= A_EXT (((std_logic_vector'("0") & (pipeline_bridge_m1_dbs_rdv_counter)) + (std_logic_vector'("0") & (pipeline_bridge_m1_dbs_rdv_counter_inc))), 2);
  --pipeline_bridge_m1_rdv_inc_mux, which is an e_mux
  pipeline_bridge_m1_dbs_rdv_counter_inc <= std_logic_vector'("01");
  --master any slave rdv, which is an e_mux
  dbs_rdv_count_enable <= pipeline_bridge_m1_read_data_valid_ext_flash_s1;
  --dbs rdv counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pipeline_bridge_m1_dbs_rdv_counter <= std_logic_vector'("00");
    elsif clk'event and clk = '1' then
      if std_logic'(dbs_rdv_count_enable) = '1' then 
        pipeline_bridge_m1_dbs_rdv_counter <= pipeline_bridge_m1_next_dbs_rdv_counter;
      end if;
    end if;

  end process;

  --dbs rdv counter overflow, which is an e_assign
  dbs_rdv_counter_overflow <= pipeline_bridge_m1_dbs_rdv_counter(1) AND NOT pipeline_bridge_m1_next_dbs_rdv_counter(1);
  --vhdl renameroo for output signals
  pipeline_bridge_m1_address_to_slave <= internal_pipeline_bridge_m1_address_to_slave;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_dbs_address <= internal_pipeline_bridge_m1_dbs_address;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_latency_counter <= internal_pipeline_bridge_m1_latency_counter;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_waitrequest <= internal_pipeline_bridge_m1_waitrequest;
--synthesis translate_off
    --pipeline_bridge_m1_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_m1_address_last_time <= std_logic_vector'("0000000000000000000000000");
      elsif clk'event and clk = '1' then
        pipeline_bridge_m1_address_last_time <= pipeline_bridge_m1_address;
      end if;

    end process;

    --pipeline_bridge/m1 waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_pipeline_bridge_m1_waitrequest AND pipeline_bridge_m1_chipselect;
      end if;

    end process;

    --pipeline_bridge_m1_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line36 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pipeline_bridge_m1_address /= pipeline_bridge_m1_address_last_time))))) = '1' then 
          write(write_line36, now);
          write(write_line36, string'(": "));
          write(write_line36, string'("pipeline_bridge_m1_address did not heed wait!!!"));
          write(output, write_line36.all);
          deallocate (write_line36);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_m1_chipselect check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_m1_chipselect_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pipeline_bridge_m1_chipselect_last_time <= pipeline_bridge_m1_chipselect;
      end if;

    end process;

    --pipeline_bridge_m1_chipselect matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line37 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pipeline_bridge_m1_chipselect) /= std_logic'(pipeline_bridge_m1_chipselect_last_time)))))) = '1' then 
          write(write_line37, now);
          write(write_line37, string'(": "));
          write(write_line37, string'("pipeline_bridge_m1_chipselect did not heed wait!!!"));
          write(output, write_line37.all);
          deallocate (write_line37);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_m1_burstcount check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_m1_burstcount_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pipeline_bridge_m1_burstcount_last_time <= pipeline_bridge_m1_burstcount;
      end if;

    end process;

    --pipeline_bridge_m1_burstcount matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line38 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pipeline_bridge_m1_burstcount) /= std_logic'(pipeline_bridge_m1_burstcount_last_time)))))) = '1' then 
          write(write_line38, now);
          write(write_line38, string'(": "));
          write(write_line38, string'("pipeline_bridge_m1_burstcount did not heed wait!!!"));
          write(output, write_line38.all);
          deallocate (write_line38);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_m1_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_m1_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        pipeline_bridge_m1_byteenable_last_time <= pipeline_bridge_m1_byteenable;
      end if;

    end process;

    --pipeline_bridge_m1_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line39 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((pipeline_bridge_m1_byteenable /= pipeline_bridge_m1_byteenable_last_time))))) = '1' then 
          write(write_line39, now);
          write(write_line39, string'(": "));
          write(write_line39, string'("pipeline_bridge_m1_byteenable did not heed wait!!!"));
          write(output, write_line39.all);
          deallocate (write_line39);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_m1_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_m1_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pipeline_bridge_m1_read_last_time <= pipeline_bridge_m1_read;
      end if;

    end process;

    --pipeline_bridge_m1_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line40 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pipeline_bridge_m1_read) /= std_logic'(pipeline_bridge_m1_read_last_time)))))) = '1' then 
          write(write_line40, now);
          write(write_line40, string'(": "));
          write(write_line40, string'("pipeline_bridge_m1_read did not heed wait!!!"));
          write(output, write_line40.all);
          deallocate (write_line40);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_m1_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_m1_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        pipeline_bridge_m1_write_last_time <= pipeline_bridge_m1_write;
      end if;

    end process;

    --pipeline_bridge_m1_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line41 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(pipeline_bridge_m1_write) /= std_logic'(pipeline_bridge_m1_write_last_time)))))) = '1' then 
          write(write_line41, now);
          write(write_line41, string'(": "));
          write(write_line41, string'("pipeline_bridge_m1_write did not heed wait!!!"));
          write(output, write_line41.all);
          deallocate (write_line41);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --pipeline_bridge_m1_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        pipeline_bridge_m1_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        pipeline_bridge_m1_writedata_last_time <= pipeline_bridge_m1_writedata;
      end if;

    end process;

    --pipeline_bridge_m1_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line42 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((pipeline_bridge_m1_writedata /= pipeline_bridge_m1_writedata_last_time)))) AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect)))) = '1' then 
          write(write_line42, now);
          write(write_line42, string'(": "));
          write(write_line42, string'("pipeline_bridge_m1_writedata did not heed wait!!!"));
          write(output, write_line42.all);
          deallocate (write_line42);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pipeline_bridge_bridge_arbitrator is 
end entity pipeline_bridge_bridge_arbitrator;


architecture europa of pipeline_bridge_bridge_arbitrator is

begin


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity pll_s1_arbitrator is 
        port (
              -- inputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal pll_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pll_s1_resetrequest : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_data_valid_pll_s1 : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1 : OUT STD_LOGIC;
                 signal d1_pll_s1_end_xfer : OUT STD_LOGIC;
                 signal pll_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal pll_s1_chipselect : OUT STD_LOGIC;
                 signal pll_s1_read : OUT STD_LOGIC;
                 signal pll_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal pll_s1_reset_n : OUT STD_LOGIC;
                 signal pll_s1_resetrequest_from_sa : OUT STD_LOGIC;
                 signal pll_s1_write : OUT STD_LOGIC;
                 signal pll_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity pll_s1_arbitrator;


architecture europa of pll_s1_arbitrator is
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_arbiterlock :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_arbiterlock2 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_continuerequest :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_saved_grant_pll_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_pll_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 :  STD_LOGIC;
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 :  STD_LOGIC;
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1 :  STD_LOGIC;
                signal pll_s1_allgrants :  STD_LOGIC;
                signal pll_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal pll_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal pll_s1_any_continuerequest :  STD_LOGIC;
                signal pll_s1_arb_counter_enable :  STD_LOGIC;
                signal pll_s1_arb_share_counter :  STD_LOGIC;
                signal pll_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal pll_s1_arb_share_set_values :  STD_LOGIC;
                signal pll_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal pll_s1_begins_xfer :  STD_LOGIC;
                signal pll_s1_end_xfer :  STD_LOGIC;
                signal pll_s1_firsttransfer :  STD_LOGIC;
                signal pll_s1_grant_vector :  STD_LOGIC;
                signal pll_s1_in_a_read_cycle :  STD_LOGIC;
                signal pll_s1_in_a_write_cycle :  STD_LOGIC;
                signal pll_s1_master_qreq_vector :  STD_LOGIC;
                signal pll_s1_non_bursting_master_requests :  STD_LOGIC;
                signal pll_s1_reg_firsttransfer :  STD_LOGIC;
                signal pll_s1_slavearbiterlockenable :  STD_LOGIC;
                signal pll_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal pll_s1_unreg_firsttransfer :  STD_LOGIC;
                signal pll_s1_waits_for_read :  STD_LOGIC;
                signal pll_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_pll_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT pll_s1_end_xfer;
    end if;

  end process;

  pll_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1);
  --assign pll_s1_readdata_from_sa = pll_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  pll_s1_readdata_from_sa <= pll_s1_readdata;
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read OR NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write)))))));
  --pll_s1_arb_share_counter set values, which is an e_mux
  pll_s1_arb_share_set_values <= std_logic'('1');
  --pll_s1_non_bursting_master_requests mux, which is an e_mux
  pll_s1_non_bursting_master_requests <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1;
  --pll_s1_any_bursting_master_saved_grant mux, which is an e_mux
  pll_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --pll_s1_arb_share_counter_next_value assignment, which is an e_assign
  pll_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(pll_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pll_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(pll_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pll_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --pll_s1_allgrants all slave grants, which is an e_mux
  pll_s1_allgrants <= pll_s1_grant_vector;
  --pll_s1_end_xfer assignment, which is an e_assign
  pll_s1_end_xfer <= NOT ((pll_s1_waits_for_read OR pll_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_pll_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_pll_s1 <= pll_s1_end_xfer AND (((NOT pll_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --pll_s1_arb_share_counter arbitration counter enable, which is an e_assign
  pll_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_pll_s1 AND pll_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_pll_s1 AND NOT pll_s1_non_bursting_master_requests));
  --pll_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pll_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(pll_s1_arb_counter_enable) = '1' then 
        pll_s1_arb_share_counter <= pll_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --pll_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pll_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((pll_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_pll_s1)) OR ((end_xfer_arb_share_counter_term_pll_s1 AND NOT pll_s1_non_bursting_master_requests)))) = '1' then 
        pll_s1_slavearbiterlockenable <= pll_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/out pll/s1 arbiterlock, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_arbiterlock <= pll_s1_slavearbiterlockenable AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_continuerequest;
  --pll_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  pll_s1_slavearbiterlockenable2 <= pll_s1_arb_share_counter_next_value;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/out pll/s1 arbiterlock2, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_arbiterlock2 <= pll_s1_slavearbiterlockenable2 AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_continuerequest;
  --pll_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  pll_s1_any_continuerequest <= std_logic'('1');
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_continuerequest continued request, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_continuerequest <= std_logic'('1');
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1;
  --pll_s1_writedata mux, which is an e_mux
  pll_s1_writedata <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata;
  --master is always granted when requested
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0/out saved-grant pll/s1, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_saved_grant_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1;
  --allow new arb cycle for pll/s1, which is an e_assign
  pll_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  pll_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  pll_s1_master_qreq_vector <= std_logic'('1');
  --pll_s1_reset_n assignment, which is an e_assign
  pll_s1_reset_n <= reset_n;
  --assign pll_s1_resetrequest_from_sa = pll_s1_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  pll_s1_resetrequest_from_sa <= pll_s1_resetrequest;
  pll_s1_chipselect <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1;
  --pll_s1_firsttransfer first transaction, which is an e_assign
  pll_s1_firsttransfer <= A_WE_StdLogic((std_logic'(pll_s1_begins_xfer) = '1'), pll_s1_unreg_firsttransfer, pll_s1_reg_firsttransfer);
  --pll_s1_unreg_firsttransfer first transaction, which is an e_assign
  pll_s1_unreg_firsttransfer <= NOT ((pll_s1_slavearbiterlockenable AND pll_s1_any_continuerequest));
  --pll_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      pll_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(pll_s1_begins_xfer) = '1' then 
        pll_s1_reg_firsttransfer <= pll_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --pll_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  pll_s1_beginbursttransfer_internal <= pll_s1_begins_xfer;
  --pll_s1_read assignment, which is an e_mux
  pll_s1_read <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read;
  --pll_s1_write assignment, which is an e_mux
  pll_s1_write <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write;
  --pll_s1_address mux, which is an e_mux
  pll_s1_address <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_nativeaddress;
  --d1_pll_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_pll_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_pll_s1_end_xfer <= pll_s1_end_xfer;
    end if;

  end process;

  --pll_s1_waits_for_read in a cycle, which is an e_mux
  pll_s1_waits_for_read <= pll_s1_in_a_read_cycle AND pll_s1_begins_xfer;
  --pll_s1_in_a_read_cycle assignment, which is an e_assign
  pll_s1_in_a_read_cycle <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= pll_s1_in_a_read_cycle;
  --pll_s1_waits_for_write in a cycle, which is an e_mux
  pll_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pll_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --pll_s1_in_a_write_cycle assignment, which is an e_assign
  pll_s1_in_a_write_cycle <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= pll_s1_in_a_write_cycle;
  wait_for_pll_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1;
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1;
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1;
--synthesis translate_off
    --pll/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity reconfig_request_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reconfig_request_pio_s1_readdata : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal d1_reconfig_request_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_reconfig_request_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_reconfig_request_pio_s1 : OUT STD_LOGIC;
                 signal reconfig_request_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal reconfig_request_pio_s1_chipselect : OUT STD_LOGIC;
                 signal reconfig_request_pio_s1_readdata_from_sa : OUT STD_LOGIC;
                 signal reconfig_request_pio_s1_reset_n : OUT STD_LOGIC;
                 signal reconfig_request_pio_s1_write_n : OUT STD_LOGIC;
                 signal reconfig_request_pio_s1_writedata : OUT STD_LOGIC
              );
end entity reconfig_request_pio_s1_arbitrator;


architecture europa of reconfig_request_pio_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_reconfig_request_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_reconfig_request_pio_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_reconfig_request_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_reconfig_request_pio_s1 :  STD_LOGIC;
                signal reconfig_request_pio_s1_allgrants :  STD_LOGIC;
                signal reconfig_request_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal reconfig_request_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal reconfig_request_pio_s1_any_continuerequest :  STD_LOGIC;
                signal reconfig_request_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal reconfig_request_pio_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal reconfig_request_pio_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal reconfig_request_pio_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal reconfig_request_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal reconfig_request_pio_s1_begins_xfer :  STD_LOGIC;
                signal reconfig_request_pio_s1_end_xfer :  STD_LOGIC;
                signal reconfig_request_pio_s1_firsttransfer :  STD_LOGIC;
                signal reconfig_request_pio_s1_grant_vector :  STD_LOGIC;
                signal reconfig_request_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal reconfig_request_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal reconfig_request_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal reconfig_request_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal reconfig_request_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal reconfig_request_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal reconfig_request_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal reconfig_request_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal reconfig_request_pio_s1_waits_for_read :  STD_LOGIC;
                signal reconfig_request_pio_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_reconfig_request_pio_s1_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_reconfig_request_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT reconfig_request_pio_s1_end_xfer;
    end if;

  end process;

  reconfig_request_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1);
  --assign reconfig_request_pio_s1_readdata_from_sa = reconfig_request_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  reconfig_request_pio_s1_readdata_from_sa <= reconfig_request_pio_s1_readdata;
  internal_pipeline_bridge_m1_requests_reconfig_request_pio_s1 <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000000001100101000000")))) AND pipeline_bridge_m1_chipselect;
  --reconfig_request_pio_s1_arb_share_counter set values, which is an e_mux
  reconfig_request_pio_s1_arb_share_set_values <= std_logic_vector'("001");
  --reconfig_request_pio_s1_non_bursting_master_requests mux, which is an e_mux
  reconfig_request_pio_s1_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_reconfig_request_pio_s1;
  --reconfig_request_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  reconfig_request_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --reconfig_request_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  reconfig_request_pio_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(reconfig_request_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (reconfig_request_pio_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(reconfig_request_pio_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (reconfig_request_pio_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --reconfig_request_pio_s1_allgrants all slave grants, which is an e_mux
  reconfig_request_pio_s1_allgrants <= reconfig_request_pio_s1_grant_vector;
  --reconfig_request_pio_s1_end_xfer assignment, which is an e_assign
  reconfig_request_pio_s1_end_xfer <= NOT ((reconfig_request_pio_s1_waits_for_read OR reconfig_request_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_reconfig_request_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_reconfig_request_pio_s1 <= reconfig_request_pio_s1_end_xfer AND (((NOT reconfig_request_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --reconfig_request_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  reconfig_request_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_reconfig_request_pio_s1 AND reconfig_request_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_reconfig_request_pio_s1 AND NOT reconfig_request_pio_s1_non_bursting_master_requests));
  --reconfig_request_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      reconfig_request_pio_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(reconfig_request_pio_s1_arb_counter_enable) = '1' then 
        reconfig_request_pio_s1_arb_share_counter <= reconfig_request_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --reconfig_request_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      reconfig_request_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((reconfig_request_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_reconfig_request_pio_s1)) OR ((end_xfer_arb_share_counter_term_reconfig_request_pio_s1 AND NOT reconfig_request_pio_s1_non_bursting_master_requests)))) = '1' then 
        reconfig_request_pio_s1_slavearbiterlockenable <= or_reduce(reconfig_request_pio_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 reconfig_request_pio/s1 arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= reconfig_request_pio_s1_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --reconfig_request_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  reconfig_request_pio_s1_slavearbiterlockenable2 <= or_reduce(reconfig_request_pio_s1_arb_share_counter_next_value);
  --pipeline_bridge/m1 reconfig_request_pio/s1 arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= reconfig_request_pio_s1_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --reconfig_request_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  reconfig_request_pio_s1_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 <= internal_pipeline_bridge_m1_requests_reconfig_request_pio_s1 AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1, which is an e_mux
  pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1 <= (internal_pipeline_bridge_m1_granted_reconfig_request_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT reconfig_request_pio_s1_waits_for_read;
  --reconfig_request_pio_s1_writedata mux, which is an e_mux
  reconfig_request_pio_s1_writedata <= pipeline_bridge_m1_writedata(0);
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_reconfig_request_pio_s1 <= internal_pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1;
  --pipeline_bridge/m1 saved-grant reconfig_request_pio/s1, which is an e_assign
  pipeline_bridge_m1_saved_grant_reconfig_request_pio_s1 <= internal_pipeline_bridge_m1_requests_reconfig_request_pio_s1;
  --allow new arb cycle for reconfig_request_pio/s1, which is an e_assign
  reconfig_request_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  reconfig_request_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  reconfig_request_pio_s1_master_qreq_vector <= std_logic'('1');
  --reconfig_request_pio_s1_reset_n assignment, which is an e_assign
  reconfig_request_pio_s1_reset_n <= reset_n;
  reconfig_request_pio_s1_chipselect <= internal_pipeline_bridge_m1_granted_reconfig_request_pio_s1;
  --reconfig_request_pio_s1_firsttransfer first transaction, which is an e_assign
  reconfig_request_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(reconfig_request_pio_s1_begins_xfer) = '1'), reconfig_request_pio_s1_unreg_firsttransfer, reconfig_request_pio_s1_reg_firsttransfer);
  --reconfig_request_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  reconfig_request_pio_s1_unreg_firsttransfer <= NOT ((reconfig_request_pio_s1_slavearbiterlockenable AND reconfig_request_pio_s1_any_continuerequest));
  --reconfig_request_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      reconfig_request_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(reconfig_request_pio_s1_begins_xfer) = '1' then 
        reconfig_request_pio_s1_reg_firsttransfer <= reconfig_request_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --reconfig_request_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  reconfig_request_pio_s1_beginbursttransfer_internal <= reconfig_request_pio_s1_begins_xfer;
  --~reconfig_request_pio_s1_write_n assignment, which is an e_mux
  reconfig_request_pio_s1_write_n <= NOT ((internal_pipeline_bridge_m1_granted_reconfig_request_pio_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect))));
  shifted_address_to_reconfig_request_pio_s1_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --reconfig_request_pio_s1_address mux, which is an e_mux
  reconfig_request_pio_s1_address <= A_EXT (A_SRL(shifted_address_to_reconfig_request_pio_s1_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_reconfig_request_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reconfig_request_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_reconfig_request_pio_s1_end_xfer <= reconfig_request_pio_s1_end_xfer;
    end if;

  end process;

  --reconfig_request_pio_s1_waits_for_read in a cycle, which is an e_mux
  reconfig_request_pio_s1_waits_for_read <= reconfig_request_pio_s1_in_a_read_cycle AND reconfig_request_pio_s1_begins_xfer;
  --reconfig_request_pio_s1_in_a_read_cycle assignment, which is an e_assign
  reconfig_request_pio_s1_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_reconfig_request_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= reconfig_request_pio_s1_in_a_read_cycle;
  --reconfig_request_pio_s1_waits_for_write in a cycle, which is an e_mux
  reconfig_request_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(reconfig_request_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --reconfig_request_pio_s1_in_a_write_cycle assignment, which is an e_assign
  reconfig_request_pio_s1_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_reconfig_request_pio_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= reconfig_request_pio_s1_in_a_write_cycle;
  wait_for_reconfig_request_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_reconfig_request_pio_s1 <= internal_pipeline_bridge_m1_granted_reconfig_request_pio_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 <= internal_pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_reconfig_request_pio_s1 <= internal_pipeline_bridge_m1_requests_reconfig_request_pio_s1;
--synthesis translate_off
    --reconfig_request_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line43 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_reconfig_request_pio_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line43, now);
          write(write_line43, string'(": "));
          write(write_line43, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave reconfig_request_pio/s1"));
          write(output, write_line43.all);
          deallocate (write_line43);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity seven_seg_pio_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal seven_seg_pio_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal d1_seven_seg_pio_s1_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_seven_seg_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_seven_seg_pio_s1 : OUT STD_LOGIC;
                 signal seven_seg_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal seven_seg_pio_s1_chipselect : OUT STD_LOGIC;
                 signal seven_seg_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal seven_seg_pio_s1_reset_n : OUT STD_LOGIC;
                 signal seven_seg_pio_s1_write_n : OUT STD_LOGIC;
                 signal seven_seg_pio_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity seven_seg_pio_s1_arbitrator;


architecture europa of seven_seg_pio_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_seven_seg_pio_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_seven_seg_pio_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_seven_seg_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_seven_seg_pio_s1 :  STD_LOGIC;
                signal seven_seg_pio_s1_allgrants :  STD_LOGIC;
                signal seven_seg_pio_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal seven_seg_pio_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal seven_seg_pio_s1_any_continuerequest :  STD_LOGIC;
                signal seven_seg_pio_s1_arb_counter_enable :  STD_LOGIC;
                signal seven_seg_pio_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal seven_seg_pio_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal seven_seg_pio_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal seven_seg_pio_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal seven_seg_pio_s1_begins_xfer :  STD_LOGIC;
                signal seven_seg_pio_s1_end_xfer :  STD_LOGIC;
                signal seven_seg_pio_s1_firsttransfer :  STD_LOGIC;
                signal seven_seg_pio_s1_grant_vector :  STD_LOGIC;
                signal seven_seg_pio_s1_in_a_read_cycle :  STD_LOGIC;
                signal seven_seg_pio_s1_in_a_write_cycle :  STD_LOGIC;
                signal seven_seg_pio_s1_master_qreq_vector :  STD_LOGIC;
                signal seven_seg_pio_s1_non_bursting_master_requests :  STD_LOGIC;
                signal seven_seg_pio_s1_reg_firsttransfer :  STD_LOGIC;
                signal seven_seg_pio_s1_slavearbiterlockenable :  STD_LOGIC;
                signal seven_seg_pio_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal seven_seg_pio_s1_unreg_firsttransfer :  STD_LOGIC;
                signal seven_seg_pio_s1_waits_for_read :  STD_LOGIC;
                signal seven_seg_pio_s1_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_seven_seg_pio_s1_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_seven_seg_pio_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT seven_seg_pio_s1_end_xfer;
    end if;

  end process;

  seven_seg_pio_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_seven_seg_pio_s1);
  --assign seven_seg_pio_s1_readdata_from_sa = seven_seg_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  seven_seg_pio_s1_readdata_from_sa <= seven_seg_pio_s1_readdata;
  internal_pipeline_bridge_m1_requests_seven_seg_pio_s1 <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 4) & std_logic_vector'("0000")) = std_logic_vector'("1000000000001000010110000")))) AND pipeline_bridge_m1_chipselect;
  --seven_seg_pio_s1_arb_share_counter set values, which is an e_mux
  seven_seg_pio_s1_arb_share_set_values <= std_logic_vector'("001");
  --seven_seg_pio_s1_non_bursting_master_requests mux, which is an e_mux
  seven_seg_pio_s1_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_seven_seg_pio_s1;
  --seven_seg_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  seven_seg_pio_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --seven_seg_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  seven_seg_pio_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(seven_seg_pio_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (seven_seg_pio_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(seven_seg_pio_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (seven_seg_pio_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --seven_seg_pio_s1_allgrants all slave grants, which is an e_mux
  seven_seg_pio_s1_allgrants <= seven_seg_pio_s1_grant_vector;
  --seven_seg_pio_s1_end_xfer assignment, which is an e_assign
  seven_seg_pio_s1_end_xfer <= NOT ((seven_seg_pio_s1_waits_for_read OR seven_seg_pio_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_seven_seg_pio_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_seven_seg_pio_s1 <= seven_seg_pio_s1_end_xfer AND (((NOT seven_seg_pio_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --seven_seg_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  seven_seg_pio_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_seven_seg_pio_s1 AND seven_seg_pio_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_seven_seg_pio_s1 AND NOT seven_seg_pio_s1_non_bursting_master_requests));
  --seven_seg_pio_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      seven_seg_pio_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(seven_seg_pio_s1_arb_counter_enable) = '1' then 
        seven_seg_pio_s1_arb_share_counter <= seven_seg_pio_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --seven_seg_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      seven_seg_pio_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((seven_seg_pio_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_seven_seg_pio_s1)) OR ((end_xfer_arb_share_counter_term_seven_seg_pio_s1 AND NOT seven_seg_pio_s1_non_bursting_master_requests)))) = '1' then 
        seven_seg_pio_s1_slavearbiterlockenable <= or_reduce(seven_seg_pio_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 seven_seg_pio/s1 arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= seven_seg_pio_s1_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --seven_seg_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  seven_seg_pio_s1_slavearbiterlockenable2 <= or_reduce(seven_seg_pio_s1_arb_share_counter_next_value);
  --pipeline_bridge/m1 seven_seg_pio/s1 arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= seven_seg_pio_s1_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --seven_seg_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  seven_seg_pio_s1_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 <= internal_pipeline_bridge_m1_requests_seven_seg_pio_s1 AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1, which is an e_mux
  pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1 <= (internal_pipeline_bridge_m1_granted_seven_seg_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT seven_seg_pio_s1_waits_for_read;
  --seven_seg_pio_s1_writedata mux, which is an e_mux
  seven_seg_pio_s1_writedata <= pipeline_bridge_m1_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_seven_seg_pio_s1 <= internal_pipeline_bridge_m1_qualified_request_seven_seg_pio_s1;
  --pipeline_bridge/m1 saved-grant seven_seg_pio/s1, which is an e_assign
  pipeline_bridge_m1_saved_grant_seven_seg_pio_s1 <= internal_pipeline_bridge_m1_requests_seven_seg_pio_s1;
  --allow new arb cycle for seven_seg_pio/s1, which is an e_assign
  seven_seg_pio_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  seven_seg_pio_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  seven_seg_pio_s1_master_qreq_vector <= std_logic'('1');
  --seven_seg_pio_s1_reset_n assignment, which is an e_assign
  seven_seg_pio_s1_reset_n <= reset_n;
  seven_seg_pio_s1_chipselect <= internal_pipeline_bridge_m1_granted_seven_seg_pio_s1;
  --seven_seg_pio_s1_firsttransfer first transaction, which is an e_assign
  seven_seg_pio_s1_firsttransfer <= A_WE_StdLogic((std_logic'(seven_seg_pio_s1_begins_xfer) = '1'), seven_seg_pio_s1_unreg_firsttransfer, seven_seg_pio_s1_reg_firsttransfer);
  --seven_seg_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  seven_seg_pio_s1_unreg_firsttransfer <= NOT ((seven_seg_pio_s1_slavearbiterlockenable AND seven_seg_pio_s1_any_continuerequest));
  --seven_seg_pio_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      seven_seg_pio_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(seven_seg_pio_s1_begins_xfer) = '1' then 
        seven_seg_pio_s1_reg_firsttransfer <= seven_seg_pio_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --seven_seg_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  seven_seg_pio_s1_beginbursttransfer_internal <= seven_seg_pio_s1_begins_xfer;
  --~seven_seg_pio_s1_write_n assignment, which is an e_mux
  seven_seg_pio_s1_write_n <= NOT ((internal_pipeline_bridge_m1_granted_seven_seg_pio_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect))));
  shifted_address_to_seven_seg_pio_s1_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --seven_seg_pio_s1_address mux, which is an e_mux
  seven_seg_pio_s1_address <= A_EXT (A_SRL(shifted_address_to_seven_seg_pio_s1_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 2);
  --d1_seven_seg_pio_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_seven_seg_pio_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_seven_seg_pio_s1_end_xfer <= seven_seg_pio_s1_end_xfer;
    end if;

  end process;

  --seven_seg_pio_s1_waits_for_read in a cycle, which is an e_mux
  seven_seg_pio_s1_waits_for_read <= seven_seg_pio_s1_in_a_read_cycle AND seven_seg_pio_s1_begins_xfer;
  --seven_seg_pio_s1_in_a_read_cycle assignment, which is an e_assign
  seven_seg_pio_s1_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_seven_seg_pio_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= seven_seg_pio_s1_in_a_read_cycle;
  --seven_seg_pio_s1_waits_for_write in a cycle, which is an e_mux
  seven_seg_pio_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(seven_seg_pio_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --seven_seg_pio_s1_in_a_write_cycle assignment, which is an e_assign
  seven_seg_pio_s1_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_seven_seg_pio_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= seven_seg_pio_s1_in_a_write_cycle;
  wait_for_seven_seg_pio_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_seven_seg_pio_s1 <= internal_pipeline_bridge_m1_granted_seven_seg_pio_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 <= internal_pipeline_bridge_m1_qualified_request_seven_seg_pio_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_seven_seg_pio_s1 <= internal_pipeline_bridge_m1_requests_seven_seg_pio_s1;
--synthesis translate_off
    --seven_seg_pio/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line44 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_seven_seg_pio_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line44, now);
          write(write_line44, string'(": "));
          write(write_line44, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave seven_seg_pio/s1"));
          write(output, write_line44.all);
          deallocate (write_line44);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_rx_csr_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_csr_irq : IN STD_LOGIC;
                 signal sgdma_rx_csr_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal d1_sgdma_rx_csr_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_sgdma_rx_csr : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_sgdma_rx_csr : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_sgdma_rx_csr : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_sgdma_rx_csr : OUT STD_LOGIC;
                 signal sgdma_rx_csr_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal sgdma_rx_csr_chipselect : OUT STD_LOGIC;
                 signal sgdma_rx_csr_irq_from_sa : OUT STD_LOGIC;
                 signal sgdma_rx_csr_read : OUT STD_LOGIC;
                 signal sgdma_rx_csr_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_csr_reset_n : OUT STD_LOGIC;
                 signal sgdma_rx_csr_write : OUT STD_LOGIC;
                 signal sgdma_rx_csr_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity sgdma_rx_csr_arbitrator;


architecture europa of sgdma_rx_csr_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sgdma_rx_csr :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_sgdma_rx_csr :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_sgdma_rx_csr :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_sgdma_rx_csr :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_sgdma_rx_csr :  STD_LOGIC;
                signal sgdma_rx_csr_allgrants :  STD_LOGIC;
                signal sgdma_rx_csr_allow_new_arb_cycle :  STD_LOGIC;
                signal sgdma_rx_csr_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sgdma_rx_csr_any_continuerequest :  STD_LOGIC;
                signal sgdma_rx_csr_arb_counter_enable :  STD_LOGIC;
                signal sgdma_rx_csr_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sgdma_rx_csr_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sgdma_rx_csr_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sgdma_rx_csr_beginbursttransfer_internal :  STD_LOGIC;
                signal sgdma_rx_csr_begins_xfer :  STD_LOGIC;
                signal sgdma_rx_csr_end_xfer :  STD_LOGIC;
                signal sgdma_rx_csr_firsttransfer :  STD_LOGIC;
                signal sgdma_rx_csr_grant_vector :  STD_LOGIC;
                signal sgdma_rx_csr_in_a_read_cycle :  STD_LOGIC;
                signal sgdma_rx_csr_in_a_write_cycle :  STD_LOGIC;
                signal sgdma_rx_csr_master_qreq_vector :  STD_LOGIC;
                signal sgdma_rx_csr_non_bursting_master_requests :  STD_LOGIC;
                signal sgdma_rx_csr_reg_firsttransfer :  STD_LOGIC;
                signal sgdma_rx_csr_slavearbiterlockenable :  STD_LOGIC;
                signal sgdma_rx_csr_slavearbiterlockenable2 :  STD_LOGIC;
                signal sgdma_rx_csr_unreg_firsttransfer :  STD_LOGIC;
                signal sgdma_rx_csr_waits_for_read :  STD_LOGIC;
                signal sgdma_rx_csr_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_sgdma_rx_csr_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_sgdma_rx_csr_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sgdma_rx_csr_end_xfer;
    end if;

  end process;

  sgdma_rx_csr_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_sgdma_rx_csr);
  --assign sgdma_rx_csr_readdata_from_sa = sgdma_rx_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sgdma_rx_csr_readdata_from_sa <= sgdma_rx_csr_readdata;
  internal_pipeline_bridge_m1_requests_sgdma_rx_csr <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 10) & std_logic_vector'("0000000000")) = std_logic_vector'("1000000000000110000000000")))) AND pipeline_bridge_m1_chipselect;
  --sgdma_rx_csr_arb_share_counter set values, which is an e_mux
  sgdma_rx_csr_arb_share_set_values <= std_logic_vector'("001");
  --sgdma_rx_csr_non_bursting_master_requests mux, which is an e_mux
  sgdma_rx_csr_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_sgdma_rx_csr;
  --sgdma_rx_csr_any_bursting_master_saved_grant mux, which is an e_mux
  sgdma_rx_csr_any_bursting_master_saved_grant <= std_logic'('0');
  --sgdma_rx_csr_arb_share_counter_next_value assignment, which is an e_assign
  sgdma_rx_csr_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sgdma_rx_csr_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sgdma_rx_csr_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sgdma_rx_csr_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sgdma_rx_csr_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --sgdma_rx_csr_allgrants all slave grants, which is an e_mux
  sgdma_rx_csr_allgrants <= sgdma_rx_csr_grant_vector;
  --sgdma_rx_csr_end_xfer assignment, which is an e_assign
  sgdma_rx_csr_end_xfer <= NOT ((sgdma_rx_csr_waits_for_read OR sgdma_rx_csr_waits_for_write));
  --end_xfer_arb_share_counter_term_sgdma_rx_csr arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sgdma_rx_csr <= sgdma_rx_csr_end_xfer AND (((NOT sgdma_rx_csr_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sgdma_rx_csr_arb_share_counter arbitration counter enable, which is an e_assign
  sgdma_rx_csr_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sgdma_rx_csr AND sgdma_rx_csr_allgrants)) OR ((end_xfer_arb_share_counter_term_sgdma_rx_csr AND NOT sgdma_rx_csr_non_bursting_master_requests));
  --sgdma_rx_csr_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_rx_csr_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(sgdma_rx_csr_arb_counter_enable) = '1' then 
        sgdma_rx_csr_arb_share_counter <= sgdma_rx_csr_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sgdma_rx_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_rx_csr_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sgdma_rx_csr_master_qreq_vector AND end_xfer_arb_share_counter_term_sgdma_rx_csr)) OR ((end_xfer_arb_share_counter_term_sgdma_rx_csr AND NOT sgdma_rx_csr_non_bursting_master_requests)))) = '1' then 
        sgdma_rx_csr_slavearbiterlockenable <= or_reduce(sgdma_rx_csr_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 sgdma_rx/csr arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= sgdma_rx_csr_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --sgdma_rx_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sgdma_rx_csr_slavearbiterlockenable2 <= or_reduce(sgdma_rx_csr_arb_share_counter_next_value);
  --pipeline_bridge/m1 sgdma_rx/csr arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= sgdma_rx_csr_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --sgdma_rx_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  sgdma_rx_csr_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_sgdma_rx_csr <= internal_pipeline_bridge_m1_requests_sgdma_rx_csr AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_sgdma_rx_csr, which is an e_mux
  pipeline_bridge_m1_read_data_valid_sgdma_rx_csr <= (internal_pipeline_bridge_m1_granted_sgdma_rx_csr AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT sgdma_rx_csr_waits_for_read;
  --sgdma_rx_csr_writedata mux, which is an e_mux
  sgdma_rx_csr_writedata <= pipeline_bridge_m1_writedata;
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_sgdma_rx_csr <= internal_pipeline_bridge_m1_qualified_request_sgdma_rx_csr;
  --pipeline_bridge/m1 saved-grant sgdma_rx/csr, which is an e_assign
  pipeline_bridge_m1_saved_grant_sgdma_rx_csr <= internal_pipeline_bridge_m1_requests_sgdma_rx_csr;
  --allow new arb cycle for sgdma_rx/csr, which is an e_assign
  sgdma_rx_csr_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sgdma_rx_csr_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sgdma_rx_csr_master_qreq_vector <= std_logic'('1');
  --sgdma_rx_csr_reset_n assignment, which is an e_assign
  sgdma_rx_csr_reset_n <= reset_n;
  sgdma_rx_csr_chipselect <= internal_pipeline_bridge_m1_granted_sgdma_rx_csr;
  --sgdma_rx_csr_firsttransfer first transaction, which is an e_assign
  sgdma_rx_csr_firsttransfer <= A_WE_StdLogic((std_logic'(sgdma_rx_csr_begins_xfer) = '1'), sgdma_rx_csr_unreg_firsttransfer, sgdma_rx_csr_reg_firsttransfer);
  --sgdma_rx_csr_unreg_firsttransfer first transaction, which is an e_assign
  sgdma_rx_csr_unreg_firsttransfer <= NOT ((sgdma_rx_csr_slavearbiterlockenable AND sgdma_rx_csr_any_continuerequest));
  --sgdma_rx_csr_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_rx_csr_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sgdma_rx_csr_begins_xfer) = '1' then 
        sgdma_rx_csr_reg_firsttransfer <= sgdma_rx_csr_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sgdma_rx_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sgdma_rx_csr_beginbursttransfer_internal <= sgdma_rx_csr_begins_xfer;
  --sgdma_rx_csr_read assignment, which is an e_mux
  sgdma_rx_csr_read <= internal_pipeline_bridge_m1_granted_sgdma_rx_csr AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --sgdma_rx_csr_write assignment, which is an e_mux
  sgdma_rx_csr_write <= internal_pipeline_bridge_m1_granted_sgdma_rx_csr AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  shifted_address_to_sgdma_rx_csr_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --sgdma_rx_csr_address mux, which is an e_mux
  sgdma_rx_csr_address <= A_EXT (A_SRL(shifted_address_to_sgdma_rx_csr_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 8);
  --d1_sgdma_rx_csr_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sgdma_rx_csr_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sgdma_rx_csr_end_xfer <= sgdma_rx_csr_end_xfer;
    end if;

  end process;

  --sgdma_rx_csr_waits_for_read in a cycle, which is an e_mux
  sgdma_rx_csr_waits_for_read <= sgdma_rx_csr_in_a_read_cycle AND sgdma_rx_csr_begins_xfer;
  --sgdma_rx_csr_in_a_read_cycle assignment, which is an e_assign
  sgdma_rx_csr_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_sgdma_rx_csr AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sgdma_rx_csr_in_a_read_cycle;
  --sgdma_rx_csr_waits_for_write in a cycle, which is an e_mux
  sgdma_rx_csr_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_rx_csr_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sgdma_rx_csr_in_a_write_cycle assignment, which is an e_assign
  sgdma_rx_csr_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_sgdma_rx_csr AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sgdma_rx_csr_in_a_write_cycle;
  wait_for_sgdma_rx_csr_counter <= std_logic'('0');
  --assign sgdma_rx_csr_irq_from_sa = sgdma_rx_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sgdma_rx_csr_irq_from_sa <= sgdma_rx_csr_irq;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_sgdma_rx_csr <= internal_pipeline_bridge_m1_granted_sgdma_rx_csr;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_sgdma_rx_csr <= internal_pipeline_bridge_m1_qualified_request_sgdma_rx_csr;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_sgdma_rx_csr <= internal_pipeline_bridge_m1_requests_sgdma_rx_csr;
--synthesis translate_off
    --sgdma_rx/csr enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line45 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_sgdma_rx_csr AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line45, now);
          write(write_line45, string'(": "));
          write(write_line45, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave sgdma_rx/csr"));
          write(output, write_line45.all);
          deallocate (write_line45);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sgdma_rx_in_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_in_ready : IN STD_LOGIC;
                 signal tse_mac_receive_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_receive_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal tse_mac_receive_endofpacket : IN STD_LOGIC;
                 signal tse_mac_receive_error : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal tse_mac_receive_startofpacket : IN STD_LOGIC;
                 signal tse_mac_receive_valid : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_rx_in_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_in_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sgdma_rx_in_endofpacket : OUT STD_LOGIC;
                 signal sgdma_rx_in_error : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal sgdma_rx_in_ready_from_sa : OUT STD_LOGIC;
                 signal sgdma_rx_in_startofpacket : OUT STD_LOGIC;
                 signal sgdma_rx_in_valid : OUT STD_LOGIC
              );
end entity sgdma_rx_in_arbitrator;


architecture europa of sgdma_rx_in_arbitrator is

begin

  --mux sgdma_rx_in_data, which is an e_mux
  sgdma_rx_in_data <= tse_mac_receive_data;
  --mux sgdma_rx_in_empty, which is an e_mux
  sgdma_rx_in_empty <= tse_mac_receive_empty;
  --mux sgdma_rx_in_endofpacket, which is an e_mux
  sgdma_rx_in_endofpacket <= tse_mac_receive_endofpacket;
  --mux sgdma_rx_in_error, which is an e_mux
  sgdma_rx_in_error <= tse_mac_receive_error;
  --assign sgdma_rx_in_ready_from_sa = sgdma_rx_in_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  sgdma_rx_in_ready_from_sa <= sgdma_rx_in_ready;
  --mux sgdma_rx_in_startofpacket, which is an e_mux
  sgdma_rx_in_startofpacket <= tse_mac_receive_startofpacket;
  --mux sgdma_rx_in_valid, which is an e_mux
  sgdma_rx_in_valid <= tse_mac_receive_valid;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_rx_descriptor_read_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                 signal descriptor_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_read_granted_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_read : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_read_requests_descriptor_memory_s1 : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_rx_descriptor_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_read_latency_counter : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_read_readdatavalid : OUT STD_LOGIC;
                 signal sgdma_rx_descriptor_read_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_rx_descriptor_read_arbitrator;


architecture europa of sgdma_rx_descriptor_read_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_rx_descriptor_read_latency_counter :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_read_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_sgdma_rx_descriptor_read_latency_counter :  STD_LOGIC;
                signal pre_flush_sgdma_rx_descriptor_read_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_read_is_granted_some_slave :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read_but_no_slave_selected :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read_last_time :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_run :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 OR NOT sgdma_rx_descriptor_read_requests_descriptor_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_descriptor_read_granted_descriptor_memory_s1 OR NOT sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 OR NOT (sgdma_rx_descriptor_read_read))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_rx_descriptor_read_read))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_rx_descriptor_read_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_rx_descriptor_read_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000100001000001000") & sgdma_rx_descriptor_read_address(12 DOWNTO 0));
  --sgdma_rx_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_rx_descriptor_read_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      sgdma_rx_descriptor_read_read_but_no_slave_selected <= (sgdma_rx_descriptor_read_read AND sgdma_rx_descriptor_read_run) AND NOT sgdma_rx_descriptor_read_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  sgdma_rx_descriptor_read_is_granted_some_slave <= sgdma_rx_descriptor_read_granted_descriptor_memory_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_sgdma_rx_descriptor_read_readdatavalid <= sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  sgdma_rx_descriptor_read_readdatavalid <= sgdma_rx_descriptor_read_read_but_no_slave_selected OR pre_flush_sgdma_rx_descriptor_read_readdatavalid;
  --sgdma_rx/descriptor_read readdata mux, which is an e_mux
  sgdma_rx_descriptor_read_readdata <= descriptor_memory_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_sgdma_rx_descriptor_read_waitrequest <= NOT sgdma_rx_descriptor_read_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_sgdma_rx_descriptor_read_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_sgdma_rx_descriptor_read_latency_counter <= p1_sgdma_rx_descriptor_read_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_sgdma_rx_descriptor_read_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((sgdma_rx_descriptor_read_run AND sgdma_rx_descriptor_read_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_sgdma_rx_descriptor_read_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_sgdma_rx_descriptor_read_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_rx_descriptor_read_requests_descriptor_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_address_to_slave <= internal_sgdma_rx_descriptor_read_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_latency_counter <= internal_sgdma_rx_descriptor_read_latency_counter;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_read_waitrequest <= internal_sgdma_rx_descriptor_read_waitrequest;
--synthesis translate_off
    --sgdma_rx_descriptor_read_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_descriptor_read_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_rx_descriptor_read_address_last_time <= sgdma_rx_descriptor_read_address;
      end if;

    end process;

    --sgdma_rx/descriptor_read waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_rx_descriptor_read_waitrequest AND (sgdma_rx_descriptor_read_read);
      end if;

    end process;

    --sgdma_rx_descriptor_read_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line46 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_descriptor_read_address /= sgdma_rx_descriptor_read_address_last_time))))) = '1' then 
          write(write_line46, now);
          write(write_line46, string'(": "));
          write(write_line46, string'("sgdma_rx_descriptor_read_address did not heed wait!!!"));
          write(output, write_line46.all);
          deallocate (write_line46);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_descriptor_read_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_descriptor_read_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_rx_descriptor_read_read_last_time <= sgdma_rx_descriptor_read_read;
      end if;

    end process;

    --sgdma_rx_descriptor_read_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line47 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_rx_descriptor_read_read) /= std_logic'(sgdma_rx_descriptor_read_read_last_time)))))) = '1' then 
          write(write_line47, now);
          write(write_line47, string'(": "));
          write(write_line47, string'("sgdma_rx_descriptor_read_read did not heed wait!!!"));
          write(output, write_line47.all);
          deallocate (write_line47);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_rx_descriptor_write_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_write_granted_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_requests_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_write : IN STD_LOGIC;
                 signal sgdma_rx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal sgdma_rx_descriptor_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_descriptor_write_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_rx_descriptor_write_arbitrator;


architecture europa of sgdma_rx_descriptor_write_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_sgdma_rx_descriptor_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_rx_descriptor_write_waitrequest :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_write_run :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_write_last_time :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 OR NOT sgdma_rx_descriptor_write_requests_descriptor_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_descriptor_write_granted_descriptor_memory_s1 OR NOT sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 OR NOT (sgdma_rx_descriptor_write_write))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_rx_descriptor_write_write))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_rx_descriptor_write_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_rx_descriptor_write_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000100001000001000") & sgdma_rx_descriptor_write_address(12 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_sgdma_rx_descriptor_write_waitrequest <= NOT sgdma_rx_descriptor_write_run;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_write_address_to_slave <= internal_sgdma_rx_descriptor_write_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_rx_descriptor_write_waitrequest <= internal_sgdma_rx_descriptor_write_waitrequest;
--synthesis translate_off
    --sgdma_rx_descriptor_write_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_descriptor_write_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_rx_descriptor_write_address_last_time <= sgdma_rx_descriptor_write_address;
      end if;

    end process;

    --sgdma_rx/descriptor_write waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_rx_descriptor_write_waitrequest AND (sgdma_rx_descriptor_write_write);
      end if;

    end process;

    --sgdma_rx_descriptor_write_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line48 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_descriptor_write_address /= sgdma_rx_descriptor_write_address_last_time))))) = '1' then 
          write(write_line48, now);
          write(write_line48, string'(": "));
          write(write_line48, string'("sgdma_rx_descriptor_write_address did not heed wait!!!"));
          write(output, write_line48.all);
          deallocate (write_line48);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_descriptor_write_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_descriptor_write_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_rx_descriptor_write_write_last_time <= sgdma_rx_descriptor_write_write;
      end if;

    end process;

    --sgdma_rx_descriptor_write_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line49 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_rx_descriptor_write_write) /= std_logic'(sgdma_rx_descriptor_write_write_last_time)))))) = '1' then 
          write(write_line49, now);
          write(write_line49, string'(": "));
          write(write_line49, string'("sgdma_rx_descriptor_write_write did not heed wait!!!"));
          write(output, write_line49.all);
          deallocate (write_line49);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_descriptor_write_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_descriptor_write_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_rx_descriptor_write_writedata_last_time <= sgdma_rx_descriptor_write_writedata;
      end if;

    end process;

    --sgdma_rx_descriptor_write_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line50 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_descriptor_write_writedata /= sgdma_rx_descriptor_write_writedata_last_time)))) AND sgdma_rx_descriptor_write_write)) = '1' then 
          write(write_line50, now);
          write(write_line50, string'(": "));
          write(write_line50, string'("sgdma_rx_descriptor_write_writedata did not heed wait!!!"));
          write(output, write_line50.all);
          deallocate (write_line50);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_rx_m_write_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_ddr_sdram_0_s1_end_xfer : IN STD_LOGIC;
                 signal d1_ext_ssram_bus_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal d1_packet_memory_s2_end_xfer : IN STD_LOGIC;
                 signal ddr_sdram_0_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_m_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal sgdma_rx_m_write_granted_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_granted_ext_ssram_s1 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_granted_packet_memory_s2 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_qualified_request_ext_ssram_s1 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_qualified_request_packet_memory_s2 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_requests_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_requests_ext_ssram_s1 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_requests_packet_memory_s2 : IN STD_LOGIC;
                 signal sgdma_rx_m_write_write : IN STD_LOGIC;
                 signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal sgdma_rx_m_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_rx_m_write_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_rx_m_write_arbitrator;


architecture europa of sgdma_rx_m_write_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_sgdma_rx_m_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_rx_m_write_waitrequest :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal sgdma_rx_m_write_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_m_write_byteenable_last_time :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sgdma_rx_m_write_run :  STD_LOGIC;
                signal sgdma_rx_m_write_write_last_time :  STD_LOGIC;
                signal sgdma_rx_m_write_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 OR NOT sgdma_rx_m_write_requests_ddr_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_m_write_granted_ddr_sdram_0_s1 OR NOT sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 OR NOT (sgdma_rx_m_write_write))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ddr_sdram_0_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_rx_m_write_write))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_rx_m_write_run <= r_0 AND r_1;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_m_write_qualified_request_ext_ssram_s1 OR NOT sgdma_rx_m_write_requests_ext_ssram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_m_write_granted_ext_ssram_s1 OR NOT sgdma_rx_m_write_qualified_request_ext_ssram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_rx_m_write_qualified_request_ext_ssram_s1 OR NOT (sgdma_rx_m_write_write))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_rx_m_write_write))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_m_write_qualified_request_packet_memory_s2 OR NOT sgdma_rx_m_write_requests_packet_memory_s2)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_rx_m_write_granted_packet_memory_s2 OR NOT sgdma_rx_m_write_qualified_request_packet_memory_s2)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_rx_m_write_qualified_request_packet_memory_s2 OR NOT (sgdma_rx_m_write_write))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_rx_m_write_write))))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_rx_m_write_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000") & A_ToStdLogicVector(sgdma_rx_m_write_address(27)) & A_ToStdLogicVector(std_logic'('0')) & sgdma_rx_m_write_address(25 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_sgdma_rx_m_write_waitrequest <= NOT sgdma_rx_m_write_run;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_address_to_slave <= internal_sgdma_rx_m_write_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_rx_m_write_waitrequest <= internal_sgdma_rx_m_write_waitrequest;
--synthesis translate_off
    --sgdma_rx_m_write_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_m_write_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_rx_m_write_address_last_time <= sgdma_rx_m_write_address;
      end if;

    end process;

    --sgdma_rx/m_write waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_rx_m_write_waitrequest AND (sgdma_rx_m_write_write);
      end if;

    end process;

    --sgdma_rx_m_write_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line51 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_m_write_address /= sgdma_rx_m_write_address_last_time))))) = '1' then 
          write(write_line51, now);
          write(write_line51, string'(": "));
          write(write_line51, string'("sgdma_rx_m_write_address did not heed wait!!!"));
          write(output, write_line51.all);
          deallocate (write_line51);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_m_write_byteenable check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_m_write_byteenable_last_time <= std_logic_vector'("0000");
      elsif clk'event and clk = '1' then
        sgdma_rx_m_write_byteenable_last_time <= sgdma_rx_m_write_byteenable;
      end if;

    end process;

    --sgdma_rx_m_write_byteenable matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line52 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_m_write_byteenable /= sgdma_rx_m_write_byteenable_last_time))))) = '1' then 
          write(write_line52, now);
          write(write_line52, string'(": "));
          write(write_line52, string'("sgdma_rx_m_write_byteenable did not heed wait!!!"));
          write(output, write_line52.all);
          deallocate (write_line52);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_m_write_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_m_write_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_rx_m_write_write_last_time <= sgdma_rx_m_write_write;
      end if;

    end process;

    --sgdma_rx_m_write_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line53 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_rx_m_write_write) /= std_logic'(sgdma_rx_m_write_write_last_time)))))) = '1' then 
          write(write_line53, now);
          write(write_line53, string'(": "));
          write(write_line53, string'("sgdma_rx_m_write_write did not heed wait!!!"));
          write(output, write_line53.all);
          deallocate (write_line53);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_rx_m_write_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_rx_m_write_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_rx_m_write_writedata_last_time <= sgdma_rx_m_write_writedata;
      end if;

    end process;

    --sgdma_rx_m_write_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line54 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((sgdma_rx_m_write_writedata /= sgdma_rx_m_write_writedata_last_time)))) AND sgdma_rx_m_write_write)) = '1' then 
          write(write_line54, now);
          write(write_line54, string'(": "));
          write(write_line54, string'("sgdma_rx_m_write_writedata did not heed wait!!!"));
          write(output, write_line54.all);
          deallocate (write_line54);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_tx_csr_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_csr_irq : IN STD_LOGIC;
                 signal sgdma_tx_csr_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal d1_sgdma_tx_csr_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_sgdma_tx_csr : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_sgdma_tx_csr : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_sgdma_tx_csr : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_sgdma_tx_csr : OUT STD_LOGIC;
                 signal sgdma_tx_csr_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal sgdma_tx_csr_chipselect : OUT STD_LOGIC;
                 signal sgdma_tx_csr_irq_from_sa : OUT STD_LOGIC;
                 signal sgdma_tx_csr_read : OUT STD_LOGIC;
                 signal sgdma_tx_csr_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_csr_reset_n : OUT STD_LOGIC;
                 signal sgdma_tx_csr_write : OUT STD_LOGIC;
                 signal sgdma_tx_csr_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity sgdma_tx_csr_arbitrator;


architecture europa of sgdma_tx_csr_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sgdma_tx_csr :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_sgdma_tx_csr :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_sgdma_tx_csr :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_sgdma_tx_csr :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_sgdma_tx_csr :  STD_LOGIC;
                signal sgdma_tx_csr_allgrants :  STD_LOGIC;
                signal sgdma_tx_csr_allow_new_arb_cycle :  STD_LOGIC;
                signal sgdma_tx_csr_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sgdma_tx_csr_any_continuerequest :  STD_LOGIC;
                signal sgdma_tx_csr_arb_counter_enable :  STD_LOGIC;
                signal sgdma_tx_csr_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sgdma_tx_csr_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sgdma_tx_csr_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sgdma_tx_csr_beginbursttransfer_internal :  STD_LOGIC;
                signal sgdma_tx_csr_begins_xfer :  STD_LOGIC;
                signal sgdma_tx_csr_end_xfer :  STD_LOGIC;
                signal sgdma_tx_csr_firsttransfer :  STD_LOGIC;
                signal sgdma_tx_csr_grant_vector :  STD_LOGIC;
                signal sgdma_tx_csr_in_a_read_cycle :  STD_LOGIC;
                signal sgdma_tx_csr_in_a_write_cycle :  STD_LOGIC;
                signal sgdma_tx_csr_master_qreq_vector :  STD_LOGIC;
                signal sgdma_tx_csr_non_bursting_master_requests :  STD_LOGIC;
                signal sgdma_tx_csr_reg_firsttransfer :  STD_LOGIC;
                signal sgdma_tx_csr_slavearbiterlockenable :  STD_LOGIC;
                signal sgdma_tx_csr_slavearbiterlockenable2 :  STD_LOGIC;
                signal sgdma_tx_csr_unreg_firsttransfer :  STD_LOGIC;
                signal sgdma_tx_csr_waits_for_read :  STD_LOGIC;
                signal sgdma_tx_csr_waits_for_write :  STD_LOGIC;
                signal shifted_address_to_sgdma_tx_csr_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal wait_for_sgdma_tx_csr_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sgdma_tx_csr_end_xfer;
    end if;

  end process;

  sgdma_tx_csr_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_sgdma_tx_csr);
  --assign sgdma_tx_csr_readdata_from_sa = sgdma_tx_csr_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sgdma_tx_csr_readdata_from_sa <= sgdma_tx_csr_readdata;
  internal_pipeline_bridge_m1_requests_sgdma_tx_csr <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 10) & std_logic_vector'("0000000000")) = std_logic_vector'("1000000000000100000000000")))) AND pipeline_bridge_m1_chipselect;
  --sgdma_tx_csr_arb_share_counter set values, which is an e_mux
  sgdma_tx_csr_arb_share_set_values <= std_logic_vector'("001");
  --sgdma_tx_csr_non_bursting_master_requests mux, which is an e_mux
  sgdma_tx_csr_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_sgdma_tx_csr;
  --sgdma_tx_csr_any_bursting_master_saved_grant mux, which is an e_mux
  sgdma_tx_csr_any_bursting_master_saved_grant <= std_logic'('0');
  --sgdma_tx_csr_arb_share_counter_next_value assignment, which is an e_assign
  sgdma_tx_csr_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sgdma_tx_csr_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sgdma_tx_csr_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sgdma_tx_csr_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sgdma_tx_csr_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --sgdma_tx_csr_allgrants all slave grants, which is an e_mux
  sgdma_tx_csr_allgrants <= sgdma_tx_csr_grant_vector;
  --sgdma_tx_csr_end_xfer assignment, which is an e_assign
  sgdma_tx_csr_end_xfer <= NOT ((sgdma_tx_csr_waits_for_read OR sgdma_tx_csr_waits_for_write));
  --end_xfer_arb_share_counter_term_sgdma_tx_csr arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sgdma_tx_csr <= sgdma_tx_csr_end_xfer AND (((NOT sgdma_tx_csr_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sgdma_tx_csr_arb_share_counter arbitration counter enable, which is an e_assign
  sgdma_tx_csr_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sgdma_tx_csr AND sgdma_tx_csr_allgrants)) OR ((end_xfer_arb_share_counter_term_sgdma_tx_csr AND NOT sgdma_tx_csr_non_bursting_master_requests));
  --sgdma_tx_csr_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_csr_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(sgdma_tx_csr_arb_counter_enable) = '1' then 
        sgdma_tx_csr_arb_share_counter <= sgdma_tx_csr_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sgdma_tx_csr_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_csr_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sgdma_tx_csr_master_qreq_vector AND end_xfer_arb_share_counter_term_sgdma_tx_csr)) OR ((end_xfer_arb_share_counter_term_sgdma_tx_csr AND NOT sgdma_tx_csr_non_bursting_master_requests)))) = '1' then 
        sgdma_tx_csr_slavearbiterlockenable <= or_reduce(sgdma_tx_csr_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 sgdma_tx/csr arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= sgdma_tx_csr_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --sgdma_tx_csr_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sgdma_tx_csr_slavearbiterlockenable2 <= or_reduce(sgdma_tx_csr_arb_share_counter_next_value);
  --pipeline_bridge/m1 sgdma_tx/csr arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= sgdma_tx_csr_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --sgdma_tx_csr_any_continuerequest at least one master continues requesting, which is an e_assign
  sgdma_tx_csr_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_sgdma_tx_csr <= internal_pipeline_bridge_m1_requests_sgdma_tx_csr AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_sgdma_tx_csr, which is an e_mux
  pipeline_bridge_m1_read_data_valid_sgdma_tx_csr <= (internal_pipeline_bridge_m1_granted_sgdma_tx_csr AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT sgdma_tx_csr_waits_for_read;
  --sgdma_tx_csr_writedata mux, which is an e_mux
  sgdma_tx_csr_writedata <= pipeline_bridge_m1_writedata;
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_sgdma_tx_csr <= internal_pipeline_bridge_m1_qualified_request_sgdma_tx_csr;
  --pipeline_bridge/m1 saved-grant sgdma_tx/csr, which is an e_assign
  pipeline_bridge_m1_saved_grant_sgdma_tx_csr <= internal_pipeline_bridge_m1_requests_sgdma_tx_csr;
  --allow new arb cycle for sgdma_tx/csr, which is an e_assign
  sgdma_tx_csr_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sgdma_tx_csr_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sgdma_tx_csr_master_qreq_vector <= std_logic'('1');
  --sgdma_tx_csr_reset_n assignment, which is an e_assign
  sgdma_tx_csr_reset_n <= reset_n;
  sgdma_tx_csr_chipselect <= internal_pipeline_bridge_m1_granted_sgdma_tx_csr;
  --sgdma_tx_csr_firsttransfer first transaction, which is an e_assign
  sgdma_tx_csr_firsttransfer <= A_WE_StdLogic((std_logic'(sgdma_tx_csr_begins_xfer) = '1'), sgdma_tx_csr_unreg_firsttransfer, sgdma_tx_csr_reg_firsttransfer);
  --sgdma_tx_csr_unreg_firsttransfer first transaction, which is an e_assign
  sgdma_tx_csr_unreg_firsttransfer <= NOT ((sgdma_tx_csr_slavearbiterlockenable AND sgdma_tx_csr_any_continuerequest));
  --sgdma_tx_csr_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_csr_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sgdma_tx_csr_begins_xfer) = '1' then 
        sgdma_tx_csr_reg_firsttransfer <= sgdma_tx_csr_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sgdma_tx_csr_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sgdma_tx_csr_beginbursttransfer_internal <= sgdma_tx_csr_begins_xfer;
  --sgdma_tx_csr_read assignment, which is an e_mux
  sgdma_tx_csr_read <= internal_pipeline_bridge_m1_granted_sgdma_tx_csr AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --sgdma_tx_csr_write assignment, which is an e_mux
  sgdma_tx_csr_write <= internal_pipeline_bridge_m1_granted_sgdma_tx_csr AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  shifted_address_to_sgdma_tx_csr_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --sgdma_tx_csr_address mux, which is an e_mux
  sgdma_tx_csr_address <= A_EXT (A_SRL(shifted_address_to_sgdma_tx_csr_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 8);
  --d1_sgdma_tx_csr_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sgdma_tx_csr_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sgdma_tx_csr_end_xfer <= sgdma_tx_csr_end_xfer;
    end if;

  end process;

  --sgdma_tx_csr_waits_for_read in a cycle, which is an e_mux
  sgdma_tx_csr_waits_for_read <= sgdma_tx_csr_in_a_read_cycle AND sgdma_tx_csr_begins_xfer;
  --sgdma_tx_csr_in_a_read_cycle assignment, which is an e_assign
  sgdma_tx_csr_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_sgdma_tx_csr AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sgdma_tx_csr_in_a_read_cycle;
  --sgdma_tx_csr_waits_for_write in a cycle, which is an e_mux
  sgdma_tx_csr_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_tx_csr_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sgdma_tx_csr_in_a_write_cycle assignment, which is an e_assign
  sgdma_tx_csr_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_sgdma_tx_csr AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sgdma_tx_csr_in_a_write_cycle;
  wait_for_sgdma_tx_csr_counter <= std_logic'('0');
  --assign sgdma_tx_csr_irq_from_sa = sgdma_tx_csr_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sgdma_tx_csr_irq_from_sa <= sgdma_tx_csr_irq;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_sgdma_tx_csr <= internal_pipeline_bridge_m1_granted_sgdma_tx_csr;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_sgdma_tx_csr <= internal_pipeline_bridge_m1_qualified_request_sgdma_tx_csr;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_sgdma_tx_csr <= internal_pipeline_bridge_m1_requests_sgdma_tx_csr;
--synthesis translate_off
    --sgdma_tx/csr enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line55 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_sgdma_tx_csr AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line55, now);
          write(write_line55, string'(": "));
          write(write_line55, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave sgdma_tx/csr"));
          write(output, write_line55.all);
          deallocate (write_line55);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_tx_descriptor_read_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                 signal descriptor_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_read_granted_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_read : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_read_requests_descriptor_memory_s1 : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_tx_descriptor_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_read_latency_counter : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_read_readdatavalid : OUT STD_LOGIC;
                 signal sgdma_tx_descriptor_read_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_tx_descriptor_read_arbitrator;


architecture europa of sgdma_tx_descriptor_read_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_tx_descriptor_read_latency_counter :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_read_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC;
                signal p1_sgdma_tx_descriptor_read_latency_counter :  STD_LOGIC;
                signal pre_flush_sgdma_tx_descriptor_read_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_read_is_granted_some_slave :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read_but_no_slave_selected :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read_last_time :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_run :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 OR NOT sgdma_tx_descriptor_read_requests_descriptor_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_descriptor_read_granted_descriptor_memory_s1 OR NOT sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 OR NOT (sgdma_tx_descriptor_read_read))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_tx_descriptor_read_read))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_tx_descriptor_read_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_tx_descriptor_read_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000100001000001000") & sgdma_tx_descriptor_read_address(12 DOWNTO 0));
  --sgdma_tx_descriptor_read_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_descriptor_read_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      sgdma_tx_descriptor_read_read_but_no_slave_selected <= (sgdma_tx_descriptor_read_read AND sgdma_tx_descriptor_read_run) AND NOT sgdma_tx_descriptor_read_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  sgdma_tx_descriptor_read_is_granted_some_slave <= sgdma_tx_descriptor_read_granted_descriptor_memory_s1;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_sgdma_tx_descriptor_read_readdatavalid <= sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1;
  --latent slave read data valid which is not flushed, which is an e_mux
  sgdma_tx_descriptor_read_readdatavalid <= sgdma_tx_descriptor_read_read_but_no_slave_selected OR pre_flush_sgdma_tx_descriptor_read_readdatavalid;
  --sgdma_tx/descriptor_read readdata mux, which is an e_mux
  sgdma_tx_descriptor_read_readdata <= descriptor_memory_s1_readdata_from_sa;
  --actual waitrequest port, which is an e_assign
  internal_sgdma_tx_descriptor_read_waitrequest <= NOT sgdma_tx_descriptor_read_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_sgdma_tx_descriptor_read_latency_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      internal_sgdma_tx_descriptor_read_latency_counter <= p1_sgdma_tx_descriptor_read_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_sgdma_tx_descriptor_read_latency_counter <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(((sgdma_tx_descriptor_read_run AND sgdma_tx_descriptor_read_read))) = '1'), (std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(latency_load_value))), A_WE_StdLogicVector((std_logic'((internal_sgdma_tx_descriptor_read_latency_counter)) = '1'), ((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(internal_sgdma_tx_descriptor_read_latency_counter))) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))));
  --read latency load values, which is an e_mux
  latency_load_value <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sgdma_tx_descriptor_read_requests_descriptor_memory_s1))) AND std_logic_vector'("00000000000000000000000000000001")));
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_address_to_slave <= internal_sgdma_tx_descriptor_read_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_latency_counter <= internal_sgdma_tx_descriptor_read_latency_counter;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_read_waitrequest <= internal_sgdma_tx_descriptor_read_waitrequest;
--synthesis translate_off
    --sgdma_tx_descriptor_read_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_descriptor_read_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_tx_descriptor_read_address_last_time <= sgdma_tx_descriptor_read_address;
      end if;

    end process;

    --sgdma_tx/descriptor_read waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_tx_descriptor_read_waitrequest AND (sgdma_tx_descriptor_read_read);
      end if;

    end process;

    --sgdma_tx_descriptor_read_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line56 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_tx_descriptor_read_address /= sgdma_tx_descriptor_read_address_last_time))))) = '1' then 
          write(write_line56, now);
          write(write_line56, string'(": "));
          write(write_line56, string'("sgdma_tx_descriptor_read_address did not heed wait!!!"));
          write(output, write_line56.all);
          deallocate (write_line56);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_tx_descriptor_read_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_descriptor_read_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_tx_descriptor_read_read_last_time <= sgdma_tx_descriptor_read_read;
      end if;

    end process;

    --sgdma_tx_descriptor_read_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line57 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_tx_descriptor_read_read) /= std_logic'(sgdma_tx_descriptor_read_read_last_time)))))) = '1' then 
          write(write_line57, now);
          write(write_line57, string'(": "));
          write(write_line57, string'("sgdma_tx_descriptor_read_read did not heed wait!!!"));
          write(output, write_line57.all);
          deallocate (write_line57);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_tx_descriptor_write_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_write_granted_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_requests_descriptor_memory_s1 : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_write : IN STD_LOGIC;
                 signal sgdma_tx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

              -- outputs:
                 signal sgdma_tx_descriptor_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_descriptor_write_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_tx_descriptor_write_arbitrator;


architecture europa of sgdma_tx_descriptor_write_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_sgdma_tx_descriptor_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_tx_descriptor_write_waitrequest :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_write_run :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_write_last_time :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_writedata_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 OR NOT sgdma_tx_descriptor_write_requests_descriptor_memory_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_descriptor_write_granted_descriptor_memory_s1 OR NOT sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 OR NOT (sgdma_tx_descriptor_write_write))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_tx_descriptor_write_write))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_tx_descriptor_write_run <= r_0;
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_tx_descriptor_write_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000100001000001000") & sgdma_tx_descriptor_write_address(12 DOWNTO 0));
  --actual waitrequest port, which is an e_assign
  internal_sgdma_tx_descriptor_write_waitrequest <= NOT sgdma_tx_descriptor_write_run;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_write_address_to_slave <= internal_sgdma_tx_descriptor_write_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_tx_descriptor_write_waitrequest <= internal_sgdma_tx_descriptor_write_waitrequest;
--synthesis translate_off
    --sgdma_tx_descriptor_write_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_descriptor_write_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_tx_descriptor_write_address_last_time <= sgdma_tx_descriptor_write_address;
      end if;

    end process;

    --sgdma_tx/descriptor_write waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_tx_descriptor_write_waitrequest AND (sgdma_tx_descriptor_write_write);
      end if;

    end process;

    --sgdma_tx_descriptor_write_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line58 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_tx_descriptor_write_address /= sgdma_tx_descriptor_write_address_last_time))))) = '1' then 
          write(write_line58, now);
          write(write_line58, string'(": "));
          write(write_line58, string'("sgdma_tx_descriptor_write_address did not heed wait!!!"));
          write(output, write_line58.all);
          deallocate (write_line58);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_tx_descriptor_write_write check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_descriptor_write_write_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_tx_descriptor_write_write_last_time <= sgdma_tx_descriptor_write_write;
      end if;

    end process;

    --sgdma_tx_descriptor_write_write matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line59 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_tx_descriptor_write_write) /= std_logic'(sgdma_tx_descriptor_write_write_last_time)))))) = '1' then 
          write(write_line59, now);
          write(write_line59, string'(": "));
          write(write_line59, string'("sgdma_tx_descriptor_write_write did not heed wait!!!"));
          write(output, write_line59.all);
          deallocate (write_line59);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_tx_descriptor_write_writedata check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_descriptor_write_writedata_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_tx_descriptor_write_writedata_last_time <= sgdma_tx_descriptor_write_writedata;
      end if;

    end process;

    --sgdma_tx_descriptor_write_writedata matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line60 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((active_and_waiting_last_time AND to_std_logic(((sgdma_tx_descriptor_write_writedata /= sgdma_tx_descriptor_write_writedata_last_time)))) AND sgdma_tx_descriptor_write_write)) = '1' then 
          write(write_line60, now);
          write(write_line60, string'(": "));
          write(write_line60, string'("sgdma_tx_descriptor_write_writedata did not heed wait!!!"));
          write(output, write_line60.all);
          deallocate (write_line60);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sgdma_tx_m_read_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal d1_ddr_sdram_0_s1_end_xfer : IN STD_LOGIC;
                 signal d1_ext_ssram_bus_avalon_slave_end_xfer : IN STD_LOGIC;
                 signal d1_packet_memory_s2_end_xfer : IN STD_LOGIC;
                 signal ddr_sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal ddr_sdram_0_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                 signal incoming_ext_ssram_bus_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal packet_memory_s2_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_m_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_granted_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_granted_ext_ssram_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_granted_packet_memory_s2 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_qualified_request_ext_ssram_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_qualified_request_packet_memory_s2 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_ext_ssram_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_read_data_valid_packet_memory_s2 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_requests_ddr_sdram_0_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_requests_ext_ssram_s1 : IN STD_LOGIC;
                 signal sgdma_tx_m_read_requests_packet_memory_s2 : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_tx_m_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_latency_counter : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal sgdma_tx_m_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_m_read_readdatavalid : OUT STD_LOGIC;
                 signal sgdma_tx_m_read_waitrequest : OUT STD_LOGIC
              );
end entity sgdma_tx_m_read_arbitrator;


architecture europa of sgdma_tx_m_read_arbitrator is
                signal active_and_waiting_last_time :  STD_LOGIC;
                signal internal_sgdma_tx_m_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_sgdma_tx_m_read_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal internal_sgdma_tx_m_read_waitrequest :  STD_LOGIC;
                signal latency_load_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal p1_sgdma_tx_m_read_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pre_flush_sgdma_tx_m_read_readdatavalid :  STD_LOGIC;
                signal r_0 :  STD_LOGIC;
                signal r_1 :  STD_LOGIC;
                signal sgdma_tx_m_read_address_last_time :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_m_read_is_granted_some_slave :  STD_LOGIC;
                signal sgdma_tx_m_read_read_but_no_slave_selected :  STD_LOGIC;
                signal sgdma_tx_m_read_read_last_time :  STD_LOGIC;
                signal sgdma_tx_m_read_run :  STD_LOGIC;

begin

  --r_0 master_run cascaded wait assignment, which is an e_assign
  r_0 <= Vector_To_Std_Logic((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 OR NOT sgdma_tx_m_read_requests_ddr_sdram_0_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_m_read_granted_ddr_sdram_0_s1 OR NOT sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 OR NOT (sgdma_tx_m_read_read))))) OR (((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(ddr_sdram_0_s1_waitrequest_n_from_sa)))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_tx_m_read_read))))))))));
  --cascaded wait assignment, which is an e_assign
  sgdma_tx_m_read_run <= r_0 AND r_1;
  --r_1 master_run cascaded wait assignment, which is an e_assign
  r_1 <= Vector_To_Std_Logic((((((((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_m_read_qualified_request_ext_ssram_s1 OR NOT sgdma_tx_m_read_requests_ext_ssram_s1)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_m_read_granted_ext_ssram_s1 OR NOT sgdma_tx_m_read_qualified_request_ext_ssram_s1)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_tx_m_read_qualified_request_ext_ssram_s1 OR NOT (sgdma_tx_m_read_read))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_tx_m_read_read))))))))) AND std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_m_read_qualified_request_packet_memory_s2 OR NOT sgdma_tx_m_read_requests_packet_memory_s2)))))) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((sgdma_tx_m_read_granted_packet_memory_s2 OR NOT sgdma_tx_m_read_qualified_request_packet_memory_s2)))))) AND (((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((NOT sgdma_tx_m_read_qualified_request_packet_memory_s2 OR NOT (sgdma_tx_m_read_read))))) OR ((std_logic_vector'("00000000000000000000000000000001") AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR((sgdma_tx_m_read_read))))))))));
  --optimize select-logic by passing only those address bits which matter.
  internal_sgdma_tx_m_read_address_to_slave <= Std_Logic_Vector'(std_logic_vector'("0000") & A_ToStdLogicVector(sgdma_tx_m_read_address(27)) & A_ToStdLogicVector(std_logic'('0')) & sgdma_tx_m_read_address(25 DOWNTO 0));
  --sgdma_tx_m_read_read_but_no_slave_selected assignment, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sgdma_tx_m_read_read_but_no_slave_selected <= std_logic'('0');
    elsif clk'event and clk = '1' then
      sgdma_tx_m_read_read_but_no_slave_selected <= (sgdma_tx_m_read_read AND sgdma_tx_m_read_run) AND NOT sgdma_tx_m_read_is_granted_some_slave;
    end if;

  end process;

  --some slave is getting selected, which is an e_mux
  sgdma_tx_m_read_is_granted_some_slave <= (sgdma_tx_m_read_granted_ddr_sdram_0_s1 OR sgdma_tx_m_read_granted_ext_ssram_s1) OR sgdma_tx_m_read_granted_packet_memory_s2;
  --latent slave read data valids which may be flushed, which is an e_mux
  pre_flush_sgdma_tx_m_read_readdatavalid <= (sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1 OR sgdma_tx_m_read_read_data_valid_ext_ssram_s1) OR sgdma_tx_m_read_read_data_valid_packet_memory_s2;
  --latent slave read data valid which is not flushed, which is an e_mux
  sgdma_tx_m_read_readdatavalid <= ((((sgdma_tx_m_read_read_but_no_slave_selected OR pre_flush_sgdma_tx_m_read_readdatavalid) OR sgdma_tx_m_read_read_but_no_slave_selected) OR pre_flush_sgdma_tx_m_read_readdatavalid) OR sgdma_tx_m_read_read_but_no_slave_selected) OR pre_flush_sgdma_tx_m_read_readdatavalid;
  --sgdma_tx/m_read readdata mux, which is an e_mux
  sgdma_tx_m_read_readdata <= (((A_REP(NOT sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1, 32) OR ddr_sdram_0_s1_readdata_from_sa)) AND ((A_REP(NOT sgdma_tx_m_read_read_data_valid_ext_ssram_s1, 32) OR incoming_ext_ssram_bus_data))) AND ((A_REP(NOT sgdma_tx_m_read_read_data_valid_packet_memory_s2, 32) OR packet_memory_s2_readdata_from_sa));
  --actual waitrequest port, which is an e_assign
  internal_sgdma_tx_m_read_waitrequest <= NOT sgdma_tx_m_read_run;
  --latent max counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      internal_sgdma_tx_m_read_latency_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      internal_sgdma_tx_m_read_latency_counter <= p1_sgdma_tx_m_read_latency_counter;
    end if;

  end process;

  --latency counter load mux, which is an e_mux
  p1_sgdma_tx_m_read_latency_counter <= A_EXT (A_WE_StdLogicVector((std_logic'(((sgdma_tx_m_read_run AND sgdma_tx_m_read_read))) = '1'), (std_logic_vector'("000000000000000000000000000000") & (latency_load_value)), A_WE_StdLogicVector((((internal_sgdma_tx_m_read_latency_counter)) /= std_logic_vector'("000")), ((std_logic_vector'("000000000000000000000000000000") & (internal_sgdma_tx_m_read_latency_counter)) - std_logic_vector'("000000000000000000000000000000001")), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --read latency load values, which is an e_mux
  latency_load_value <= A_EXT (((((std_logic_vector'("00000000000000000000000000000") & (A_REP(sgdma_tx_m_read_requests_ext_ssram_s1, 3))) AND std_logic_vector'("00000000000000000000000000000101"))) OR (((std_logic_vector'("00000000000000000000000000000") & (A_REP(sgdma_tx_m_read_requests_packet_memory_s2, 3))) AND std_logic_vector'("00000000000000000000000000000001")))), 3);
  --vhdl renameroo for output signals
  sgdma_tx_m_read_address_to_slave <= internal_sgdma_tx_m_read_address_to_slave;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_latency_counter <= internal_sgdma_tx_m_read_latency_counter;
  --vhdl renameroo for output signals
  sgdma_tx_m_read_waitrequest <= internal_sgdma_tx_m_read_waitrequest;
--synthesis translate_off
    --sgdma_tx_m_read_address check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_m_read_address_last_time <= std_logic_vector'("00000000000000000000000000000000");
      elsif clk'event and clk = '1' then
        sgdma_tx_m_read_address_last_time <= sgdma_tx_m_read_address;
      end if;

    end process;

    --sgdma_tx/m_read waited last time, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        active_and_waiting_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        active_and_waiting_last_time <= internal_sgdma_tx_m_read_waitrequest AND (sgdma_tx_m_read_read);
      end if;

    end process;

    --sgdma_tx_m_read_address matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line61 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((sgdma_tx_m_read_address /= sgdma_tx_m_read_address_last_time))))) = '1' then 
          write(write_line61, now);
          write(write_line61, string'(": "));
          write(write_line61, string'("sgdma_tx_m_read_address did not heed wait!!!"));
          write(output, write_line61.all);
          deallocate (write_line61);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

    --sgdma_tx_m_read_read check against wait, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        sgdma_tx_m_read_read_last_time <= std_logic'('0');
      elsif clk'event and clk = '1' then
        sgdma_tx_m_read_read_last_time <= sgdma_tx_m_read_read;
      end if;

    end process;

    --sgdma_tx_m_read_read matches last port_name, which is an e_process
    process (clk)
    VARIABLE write_line62 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'((active_and_waiting_last_time AND to_std_logic(((std_logic'(sgdma_tx_m_read_read) /= std_logic'(sgdma_tx_m_read_read_last_time)))))) = '1' then 
          write(write_line62, now);
          write(write_line62, string'(": "));
          write(write_line62, string'("sgdma_tx_m_read_read did not heed wait!!!"));
          write(output, write_line62.all);
          deallocate (write_line62);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity sgdma_tx_out_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sgdma_tx_out_endofpacket : IN STD_LOGIC;
                 signal sgdma_tx_out_error : IN STD_LOGIC;
                 signal sgdma_tx_out_startofpacket : IN STD_LOGIC;
                 signal sgdma_tx_out_valid : IN STD_LOGIC;
                 signal tse_mac_transmit_ready_from_sa : IN STD_LOGIC;

              -- outputs:
                 signal sgdma_tx_out_ready : OUT STD_LOGIC
              );
end entity sgdma_tx_out_arbitrator;


architecture europa of sgdma_tx_out_arbitrator is

begin

  --mux sgdma_tx_out_ready, which is an e_mux
  sgdma_tx_out_ready <= tse_mac_transmit_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity sys_clk_timer_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal sys_clk_timer_s1_irq : IN STD_LOGIC;
                 signal sys_clk_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- outputs:
                 signal d1_sys_clk_timer_s1_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_sys_clk_timer_s1 : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal sys_clk_timer_s1_chipselect : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_irq_from_sa : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal sys_clk_timer_s1_reset_n : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_write_n : OUT STD_LOGIC;
                 signal sys_clk_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity sys_clk_timer_s1_arbitrator;


architecture europa of sys_clk_timer_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_sys_clk_timer_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_sys_clk_timer_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_sys_clk_timer_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_sys_clk_timer_s1 :  STD_LOGIC;
                signal shifted_address_to_sys_clk_timer_s1_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal sys_clk_timer_s1_allgrants :  STD_LOGIC;
                signal sys_clk_timer_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal sys_clk_timer_s1_any_continuerequest :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_counter_enable :  STD_LOGIC;
                signal sys_clk_timer_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sys_clk_timer_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sys_clk_timer_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sys_clk_timer_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal sys_clk_timer_s1_begins_xfer :  STD_LOGIC;
                signal sys_clk_timer_s1_end_xfer :  STD_LOGIC;
                signal sys_clk_timer_s1_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_grant_vector :  STD_LOGIC;
                signal sys_clk_timer_s1_in_a_read_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_in_a_write_cycle :  STD_LOGIC;
                signal sys_clk_timer_s1_master_qreq_vector :  STD_LOGIC;
                signal sys_clk_timer_s1_non_bursting_master_requests :  STD_LOGIC;
                signal sys_clk_timer_s1_reg_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_slavearbiterlockenable :  STD_LOGIC;
                signal sys_clk_timer_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal sys_clk_timer_s1_unreg_firsttransfer :  STD_LOGIC;
                signal sys_clk_timer_s1_waits_for_read :  STD_LOGIC;
                signal sys_clk_timer_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_sys_clk_timer_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT sys_clk_timer_s1_end_xfer;
    end if;

  end process;

  sys_clk_timer_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_sys_clk_timer_s1);
  --assign sys_clk_timer_s1_readdata_from_sa = sys_clk_timer_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  sys_clk_timer_s1_readdata_from_sa <= sys_clk_timer_s1_readdata;
  internal_pipeline_bridge_m1_requests_sys_clk_timer_s1 <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1000000000001000001100000")))) AND pipeline_bridge_m1_chipselect;
  --sys_clk_timer_s1_arb_share_counter set values, which is an e_mux
  sys_clk_timer_s1_arb_share_set_values <= std_logic_vector'("001");
  --sys_clk_timer_s1_non_bursting_master_requests mux, which is an e_mux
  sys_clk_timer_s1_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_sys_clk_timer_s1;
  --sys_clk_timer_s1_any_bursting_master_saved_grant mux, which is an e_mux
  sys_clk_timer_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --sys_clk_timer_s1_arb_share_counter_next_value assignment, which is an e_assign
  sys_clk_timer_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(sys_clk_timer_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sys_clk_timer_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(sys_clk_timer_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (sys_clk_timer_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --sys_clk_timer_s1_allgrants all slave grants, which is an e_mux
  sys_clk_timer_s1_allgrants <= sys_clk_timer_s1_grant_vector;
  --sys_clk_timer_s1_end_xfer assignment, which is an e_assign
  sys_clk_timer_s1_end_xfer <= NOT ((sys_clk_timer_s1_waits_for_read OR sys_clk_timer_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_sys_clk_timer_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_sys_clk_timer_s1 <= sys_clk_timer_s1_end_xfer AND (((NOT sys_clk_timer_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --sys_clk_timer_s1_arb_share_counter arbitration counter enable, which is an e_assign
  sys_clk_timer_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND sys_clk_timer_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND NOT sys_clk_timer_s1_non_bursting_master_requests));
  --sys_clk_timer_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(sys_clk_timer_s1_arb_counter_enable) = '1' then 
        sys_clk_timer_s1_arb_share_counter <= sys_clk_timer_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --sys_clk_timer_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((sys_clk_timer_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_sys_clk_timer_s1)) OR ((end_xfer_arb_share_counter_term_sys_clk_timer_s1 AND NOT sys_clk_timer_s1_non_bursting_master_requests)))) = '1' then 
        sys_clk_timer_s1_slavearbiterlockenable <= or_reduce(sys_clk_timer_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 sys_clk_timer/s1 arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= sys_clk_timer_s1_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --sys_clk_timer_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  sys_clk_timer_s1_slavearbiterlockenable2 <= or_reduce(sys_clk_timer_s1_arb_share_counter_next_value);
  --pipeline_bridge/m1 sys_clk_timer/s1 arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= sys_clk_timer_s1_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --sys_clk_timer_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  sys_clk_timer_s1_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 <= internal_pipeline_bridge_m1_requests_sys_clk_timer_s1 AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1, which is an e_mux
  pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1 <= (internal_pipeline_bridge_m1_granted_sys_clk_timer_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT sys_clk_timer_s1_waits_for_read;
  --sys_clk_timer_s1_writedata mux, which is an e_mux
  sys_clk_timer_s1_writedata <= pipeline_bridge_m1_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_sys_clk_timer_s1 <= internal_pipeline_bridge_m1_qualified_request_sys_clk_timer_s1;
  --pipeline_bridge/m1 saved-grant sys_clk_timer/s1, which is an e_assign
  pipeline_bridge_m1_saved_grant_sys_clk_timer_s1 <= internal_pipeline_bridge_m1_requests_sys_clk_timer_s1;
  --allow new arb cycle for sys_clk_timer/s1, which is an e_assign
  sys_clk_timer_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  sys_clk_timer_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  sys_clk_timer_s1_master_qreq_vector <= std_logic'('1');
  --sys_clk_timer_s1_reset_n assignment, which is an e_assign
  sys_clk_timer_s1_reset_n <= reset_n;
  sys_clk_timer_s1_chipselect <= internal_pipeline_bridge_m1_granted_sys_clk_timer_s1;
  --sys_clk_timer_s1_firsttransfer first transaction, which is an e_assign
  sys_clk_timer_s1_firsttransfer <= A_WE_StdLogic((std_logic'(sys_clk_timer_s1_begins_xfer) = '1'), sys_clk_timer_s1_unreg_firsttransfer, sys_clk_timer_s1_reg_firsttransfer);
  --sys_clk_timer_s1_unreg_firsttransfer first transaction, which is an e_assign
  sys_clk_timer_s1_unreg_firsttransfer <= NOT ((sys_clk_timer_s1_slavearbiterlockenable AND sys_clk_timer_s1_any_continuerequest));
  --sys_clk_timer_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      sys_clk_timer_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(sys_clk_timer_s1_begins_xfer) = '1' then 
        sys_clk_timer_s1_reg_firsttransfer <= sys_clk_timer_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --sys_clk_timer_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  sys_clk_timer_s1_beginbursttransfer_internal <= sys_clk_timer_s1_begins_xfer;
  --~sys_clk_timer_s1_write_n assignment, which is an e_mux
  sys_clk_timer_s1_write_n <= NOT ((internal_pipeline_bridge_m1_granted_sys_clk_timer_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect))));
  shifted_address_to_sys_clk_timer_s1_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --sys_clk_timer_s1_address mux, which is an e_mux
  sys_clk_timer_s1_address <= A_EXT (A_SRL(shifted_address_to_sys_clk_timer_s1_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_sys_clk_timer_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_sys_clk_timer_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_sys_clk_timer_s1_end_xfer <= sys_clk_timer_s1_end_xfer;
    end if;

  end process;

  --sys_clk_timer_s1_waits_for_read in a cycle, which is an e_mux
  sys_clk_timer_s1_waits_for_read <= sys_clk_timer_s1_in_a_read_cycle AND sys_clk_timer_s1_begins_xfer;
  --sys_clk_timer_s1_in_a_read_cycle assignment, which is an e_assign
  sys_clk_timer_s1_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_sys_clk_timer_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= sys_clk_timer_s1_in_a_read_cycle;
  --sys_clk_timer_s1_waits_for_write in a cycle, which is an e_mux
  sys_clk_timer_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(sys_clk_timer_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --sys_clk_timer_s1_in_a_write_cycle assignment, which is an e_assign
  sys_clk_timer_s1_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_sys_clk_timer_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= sys_clk_timer_s1_in_a_write_cycle;
  wait_for_sys_clk_timer_s1_counter <= std_logic'('0');
  --assign sys_clk_timer_s1_irq_from_sa = sys_clk_timer_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  sys_clk_timer_s1_irq_from_sa <= sys_clk_timer_s1_irq;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_sys_clk_timer_s1 <= internal_pipeline_bridge_m1_granted_sys_clk_timer_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 <= internal_pipeline_bridge_m1_qualified_request_sys_clk_timer_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_sys_clk_timer_s1 <= internal_pipeline_bridge_m1_requests_sys_clk_timer_s1;
--synthesis translate_off
    --sys_clk_timer/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line63 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_sys_clk_timer_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line63, now);
          write(write_line63, string'(": "));
          write(write_line63, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave sys_clk_timer/s1"));
          write(output, write_line63.all);
          deallocate (write_line63);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tse_mac_control_port_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                 signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal cpu_data_master_read : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                 signal cpu_data_master_write : IN STD_LOGIC;
                 signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal tse_mac_control_port_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_control_port_waitrequest : IN STD_LOGIC;

              -- outputs:
                 signal cpu_data_master_granted_tse_mac_control_port : OUT STD_LOGIC;
                 signal cpu_data_master_qualified_request_tse_mac_control_port : OUT STD_LOGIC;
                 signal cpu_data_master_read_data_valid_tse_mac_control_port : OUT STD_LOGIC;
                 signal cpu_data_master_requests_tse_mac_control_port : OUT STD_LOGIC;
                 signal d1_tse_mac_control_port_end_xfer : OUT STD_LOGIC;
                 signal tse_mac_control_port_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal tse_mac_control_port_read : OUT STD_LOGIC;
                 signal tse_mac_control_port_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_control_port_reset : OUT STD_LOGIC;
                 signal tse_mac_control_port_waitrequest_from_sa : OUT STD_LOGIC;
                 signal tse_mac_control_port_write : OUT STD_LOGIC;
                 signal tse_mac_control_port_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity tse_mac_control_port_arbitrator;


architecture europa of tse_mac_control_port_arbitrator is
                signal cpu_data_master_arbiterlock :  STD_LOGIC;
                signal cpu_data_master_arbiterlock2 :  STD_LOGIC;
                signal cpu_data_master_continuerequest :  STD_LOGIC;
                signal cpu_data_master_saved_grant_tse_mac_control_port :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_tse_mac_control_port :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_cpu_data_master_granted_tse_mac_control_port :  STD_LOGIC;
                signal internal_cpu_data_master_qualified_request_tse_mac_control_port :  STD_LOGIC;
                signal internal_cpu_data_master_requests_tse_mac_control_port :  STD_LOGIC;
                signal internal_tse_mac_control_port_waitrequest_from_sa :  STD_LOGIC;
                signal shifted_address_to_tse_mac_control_port_from_cpu_data_master :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal tse_mac_control_port_allgrants :  STD_LOGIC;
                signal tse_mac_control_port_allow_new_arb_cycle :  STD_LOGIC;
                signal tse_mac_control_port_any_bursting_master_saved_grant :  STD_LOGIC;
                signal tse_mac_control_port_any_continuerequest :  STD_LOGIC;
                signal tse_mac_control_port_arb_counter_enable :  STD_LOGIC;
                signal tse_mac_control_port_arb_share_counter :  STD_LOGIC;
                signal tse_mac_control_port_arb_share_counter_next_value :  STD_LOGIC;
                signal tse_mac_control_port_arb_share_set_values :  STD_LOGIC;
                signal tse_mac_control_port_beginbursttransfer_internal :  STD_LOGIC;
                signal tse_mac_control_port_begins_xfer :  STD_LOGIC;
                signal tse_mac_control_port_end_xfer :  STD_LOGIC;
                signal tse_mac_control_port_firsttransfer :  STD_LOGIC;
                signal tse_mac_control_port_grant_vector :  STD_LOGIC;
                signal tse_mac_control_port_in_a_read_cycle :  STD_LOGIC;
                signal tse_mac_control_port_in_a_write_cycle :  STD_LOGIC;
                signal tse_mac_control_port_master_qreq_vector :  STD_LOGIC;
                signal tse_mac_control_port_non_bursting_master_requests :  STD_LOGIC;
                signal tse_mac_control_port_reg_firsttransfer :  STD_LOGIC;
                signal tse_mac_control_port_slavearbiterlockenable :  STD_LOGIC;
                signal tse_mac_control_port_slavearbiterlockenable2 :  STD_LOGIC;
                signal tse_mac_control_port_unreg_firsttransfer :  STD_LOGIC;
                signal tse_mac_control_port_waits_for_read :  STD_LOGIC;
                signal tse_mac_control_port_waits_for_write :  STD_LOGIC;
                signal wait_for_tse_mac_control_port_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT tse_mac_control_port_end_xfer;
    end if;

  end process;

  tse_mac_control_port_begins_xfer <= NOT d1_reasons_to_wait AND (internal_cpu_data_master_qualified_request_tse_mac_control_port);
  --assign tse_mac_control_port_readdata_from_sa = tse_mac_control_port_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  tse_mac_control_port_readdata_from_sa <= tse_mac_control_port_readdata;
  internal_cpu_data_master_requests_tse_mac_control_port <= to_std_logic(((Std_Logic_Vector'(cpu_data_master_address_to_slave(27 DOWNTO 10) & std_logic_vector'("0000000000")) = std_logic_vector'("1000010000010010000000000000")))) AND ((cpu_data_master_read OR cpu_data_master_write));
  --assign tse_mac_control_port_waitrequest_from_sa = tse_mac_control_port_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  internal_tse_mac_control_port_waitrequest_from_sa <= tse_mac_control_port_waitrequest;
  --tse_mac_control_port_arb_share_counter set values, which is an e_mux
  tse_mac_control_port_arb_share_set_values <= std_logic'('1');
  --tse_mac_control_port_non_bursting_master_requests mux, which is an e_mux
  tse_mac_control_port_non_bursting_master_requests <= internal_cpu_data_master_requests_tse_mac_control_port;
  --tse_mac_control_port_any_bursting_master_saved_grant mux, which is an e_mux
  tse_mac_control_port_any_bursting_master_saved_grant <= std_logic'('0');
  --tse_mac_control_port_arb_share_counter_next_value assignment, which is an e_assign
  tse_mac_control_port_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(tse_mac_control_port_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_mac_control_port_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(tse_mac_control_port_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_mac_control_port_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --tse_mac_control_port_allgrants all slave grants, which is an e_mux
  tse_mac_control_port_allgrants <= tse_mac_control_port_grant_vector;
  --tse_mac_control_port_end_xfer assignment, which is an e_assign
  tse_mac_control_port_end_xfer <= NOT ((tse_mac_control_port_waits_for_read OR tse_mac_control_port_waits_for_write));
  --end_xfer_arb_share_counter_term_tse_mac_control_port arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_tse_mac_control_port <= tse_mac_control_port_end_xfer AND (((NOT tse_mac_control_port_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --tse_mac_control_port_arb_share_counter arbitration counter enable, which is an e_assign
  tse_mac_control_port_arb_counter_enable <= ((end_xfer_arb_share_counter_term_tse_mac_control_port AND tse_mac_control_port_allgrants)) OR ((end_xfer_arb_share_counter_term_tse_mac_control_port AND NOT tse_mac_control_port_non_bursting_master_requests));
  --tse_mac_control_port_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_mac_control_port_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(tse_mac_control_port_arb_counter_enable) = '1' then 
        tse_mac_control_port_arb_share_counter <= tse_mac_control_port_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --tse_mac_control_port_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_mac_control_port_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((tse_mac_control_port_master_qreq_vector AND end_xfer_arb_share_counter_term_tse_mac_control_port)) OR ((end_xfer_arb_share_counter_term_tse_mac_control_port AND NOT tse_mac_control_port_non_bursting_master_requests)))) = '1' then 
        tse_mac_control_port_slavearbiterlockenable <= tse_mac_control_port_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --cpu/data_master tse_mac/control_port arbiterlock, which is an e_assign
  cpu_data_master_arbiterlock <= tse_mac_control_port_slavearbiterlockenable AND cpu_data_master_continuerequest;
  --tse_mac_control_port_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  tse_mac_control_port_slavearbiterlockenable2 <= tse_mac_control_port_arb_share_counter_next_value;
  --cpu/data_master tse_mac/control_port arbiterlock2, which is an e_assign
  cpu_data_master_arbiterlock2 <= tse_mac_control_port_slavearbiterlockenable2 AND cpu_data_master_continuerequest;
  --tse_mac_control_port_any_continuerequest at least one master continues requesting, which is an e_assign
  tse_mac_control_port_any_continuerequest <= std_logic'('1');
  --cpu_data_master_continuerequest continued request, which is an e_assign
  cpu_data_master_continuerequest <= std_logic'('1');
  internal_cpu_data_master_qualified_request_tse_mac_control_port <= internal_cpu_data_master_requests_tse_mac_control_port AND NOT ((cpu_data_master_read AND (((to_std_logic((((std_logic_vector'("00000000000000000000000000000") & (cpu_data_master_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000")))) OR (cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register)) OR (cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register)))));
  --local readdatavalid cpu_data_master_read_data_valid_tse_mac_control_port, which is an e_mux
  cpu_data_master_read_data_valid_tse_mac_control_port <= (internal_cpu_data_master_granted_tse_mac_control_port AND cpu_data_master_read) AND NOT tse_mac_control_port_waits_for_read;
  --tse_mac_control_port_writedata mux, which is an e_mux
  tse_mac_control_port_writedata <= cpu_data_master_writedata;
  --master is always granted when requested
  internal_cpu_data_master_granted_tse_mac_control_port <= internal_cpu_data_master_qualified_request_tse_mac_control_port;
  --cpu/data_master saved-grant tse_mac/control_port, which is an e_assign
  cpu_data_master_saved_grant_tse_mac_control_port <= internal_cpu_data_master_requests_tse_mac_control_port;
  --allow new arb cycle for tse_mac/control_port, which is an e_assign
  tse_mac_control_port_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  tse_mac_control_port_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  tse_mac_control_port_master_qreq_vector <= std_logic'('1');
  --~tse_mac_control_port_reset assignment, which is an e_assign
  tse_mac_control_port_reset <= NOT reset_n;
  --tse_mac_control_port_firsttransfer first transaction, which is an e_assign
  tse_mac_control_port_firsttransfer <= A_WE_StdLogic((std_logic'(tse_mac_control_port_begins_xfer) = '1'), tse_mac_control_port_unreg_firsttransfer, tse_mac_control_port_reg_firsttransfer);
  --tse_mac_control_port_unreg_firsttransfer first transaction, which is an e_assign
  tse_mac_control_port_unreg_firsttransfer <= NOT ((tse_mac_control_port_slavearbiterlockenable AND tse_mac_control_port_any_continuerequest));
  --tse_mac_control_port_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_mac_control_port_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(tse_mac_control_port_begins_xfer) = '1' then 
        tse_mac_control_port_reg_firsttransfer <= tse_mac_control_port_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --tse_mac_control_port_beginbursttransfer_internal begin burst transfer, which is an e_assign
  tse_mac_control_port_beginbursttransfer_internal <= tse_mac_control_port_begins_xfer;
  --tse_mac_control_port_read assignment, which is an e_mux
  tse_mac_control_port_read <= internal_cpu_data_master_granted_tse_mac_control_port AND cpu_data_master_read;
  --tse_mac_control_port_write assignment, which is an e_mux
  tse_mac_control_port_write <= internal_cpu_data_master_granted_tse_mac_control_port AND cpu_data_master_write;
  shifted_address_to_tse_mac_control_port_from_cpu_data_master <= cpu_data_master_address_to_slave;
  --tse_mac_control_port_address mux, which is an e_mux
  tse_mac_control_port_address <= A_EXT (A_SRL(shifted_address_to_tse_mac_control_port_from_cpu_data_master,std_logic_vector'("00000000000000000000000000000010")), 8);
  --d1_tse_mac_control_port_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_tse_mac_control_port_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_tse_mac_control_port_end_xfer <= tse_mac_control_port_end_xfer;
    end if;

  end process;

  --tse_mac_control_port_waits_for_read in a cycle, which is an e_mux
  tse_mac_control_port_waits_for_read <= tse_mac_control_port_in_a_read_cycle AND internal_tse_mac_control_port_waitrequest_from_sa;
  --tse_mac_control_port_in_a_read_cycle assignment, which is an e_assign
  tse_mac_control_port_in_a_read_cycle <= internal_cpu_data_master_granted_tse_mac_control_port AND cpu_data_master_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= tse_mac_control_port_in_a_read_cycle;
  --tse_mac_control_port_waits_for_write in a cycle, which is an e_mux
  tse_mac_control_port_waits_for_write <= tse_mac_control_port_in_a_write_cycle AND internal_tse_mac_control_port_waitrequest_from_sa;
  --tse_mac_control_port_in_a_write_cycle assignment, which is an e_assign
  tse_mac_control_port_in_a_write_cycle <= internal_cpu_data_master_granted_tse_mac_control_port AND cpu_data_master_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= tse_mac_control_port_in_a_write_cycle;
  wait_for_tse_mac_control_port_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  cpu_data_master_granted_tse_mac_control_port <= internal_cpu_data_master_granted_tse_mac_control_port;
  --vhdl renameroo for output signals
  cpu_data_master_qualified_request_tse_mac_control_port <= internal_cpu_data_master_qualified_request_tse_mac_control_port;
  --vhdl renameroo for output signals
  cpu_data_master_requests_tse_mac_control_port <= internal_cpu_data_master_requests_tse_mac_control_port;
  --vhdl renameroo for output signals
  tse_mac_control_port_waitrequest_from_sa <= internal_tse_mac_control_port_waitrequest_from_sa;
--synthesis translate_off
    --tse_mac/control_port enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tse_mac_transmit_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_tx_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal sgdma_tx_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal sgdma_tx_out_endofpacket : IN STD_LOGIC;
                 signal sgdma_tx_out_error : IN STD_LOGIC;
                 signal sgdma_tx_out_startofpacket : IN STD_LOGIC;
                 signal sgdma_tx_out_valid : IN STD_LOGIC;
                 signal tse_mac_transmit_ready : IN STD_LOGIC;

              -- outputs:
                 signal tse_mac_transmit_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_transmit_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal tse_mac_transmit_endofpacket : OUT STD_LOGIC;
                 signal tse_mac_transmit_error : OUT STD_LOGIC;
                 signal tse_mac_transmit_ready_from_sa : OUT STD_LOGIC;
                 signal tse_mac_transmit_startofpacket : OUT STD_LOGIC;
                 signal tse_mac_transmit_valid : OUT STD_LOGIC
              );
end entity tse_mac_transmit_arbitrator;


architecture europa of tse_mac_transmit_arbitrator is

begin

  --mux tse_mac_transmit_data, which is an e_mux
  tse_mac_transmit_data <= sgdma_tx_out_data;
  --mux tse_mac_transmit_endofpacket, which is an e_mux
  tse_mac_transmit_endofpacket <= sgdma_tx_out_endofpacket;
  --mux tse_mac_transmit_error, which is an e_mux
  tse_mac_transmit_error <= sgdma_tx_out_error;
  --mux tse_mac_transmit_empty, which is an e_mux
  tse_mac_transmit_empty <= sgdma_tx_out_empty;
  --assign tse_mac_transmit_ready_from_sa = tse_mac_transmit_ready so that symbol knows where to group signals which may go to master only, which is an e_assign
  tse_mac_transmit_ready_from_sa <= tse_mac_transmit_ready;
  --mux tse_mac_transmit_startofpacket, which is an e_mux
  tse_mac_transmit_startofpacket <= sgdma_tx_out_startofpacket;
  --mux tse_mac_transmit_valid, which is an e_mux
  tse_mac_transmit_valid <= sgdma_tx_out_valid;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tse_mac_receive_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal sgdma_rx_in_ready_from_sa : IN STD_LOGIC;
                 signal tse_mac_receive_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal tse_mac_receive_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal tse_mac_receive_endofpacket : IN STD_LOGIC;
                 signal tse_mac_receive_error : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal tse_mac_receive_startofpacket : IN STD_LOGIC;
                 signal tse_mac_receive_valid : IN STD_LOGIC;

              -- outputs:
                 signal tse_mac_receive_ready : OUT STD_LOGIC
              );
end entity tse_mac_receive_arbitrator;


architecture europa of tse_mac_receive_arbitrator is

begin

  --mux tse_mac_receive_ready, which is an e_mux
  tse_mac_receive_ready <= sgdma_rx_in_ready_from_sa;

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity tse_pll_s1_arbitrator is 
        port (
              -- inputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write : IN STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal clk : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal tse_pll_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal tse_pll_s1_resetrequest : IN STD_LOGIC;

              -- outputs:
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_data_valid_tse_pll_s1 : OUT STD_LOGIC;
                 signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1 : OUT STD_LOGIC;
                 signal d1_tse_pll_s1_end_xfer : OUT STD_LOGIC;
                 signal tse_pll_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal tse_pll_s1_chipselect : OUT STD_LOGIC;
                 signal tse_pll_s1_read : OUT STD_LOGIC;
                 signal tse_pll_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal tse_pll_s1_reset_n : OUT STD_LOGIC;
                 signal tse_pll_s1_resetrequest_from_sa : OUT STD_LOGIC;
                 signal tse_pll_s1_write : OUT STD_LOGIC;
                 signal tse_pll_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity tse_pll_s1_arbitrator;


architecture europa of tse_pll_s1_arbitrator is
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_arbiterlock :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_arbiterlock2 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_continuerequest :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_saved_grant_tse_pll_s1 :  STD_LOGIC;
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_tse_pll_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 :  STD_LOGIC;
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 :  STD_LOGIC;
                signal internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1 :  STD_LOGIC;
                signal tse_pll_s1_allgrants :  STD_LOGIC;
                signal tse_pll_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal tse_pll_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal tse_pll_s1_any_continuerequest :  STD_LOGIC;
                signal tse_pll_s1_arb_counter_enable :  STD_LOGIC;
                signal tse_pll_s1_arb_share_counter :  STD_LOGIC;
                signal tse_pll_s1_arb_share_counter_next_value :  STD_LOGIC;
                signal tse_pll_s1_arb_share_set_values :  STD_LOGIC;
                signal tse_pll_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal tse_pll_s1_begins_xfer :  STD_LOGIC;
                signal tse_pll_s1_end_xfer :  STD_LOGIC;
                signal tse_pll_s1_firsttransfer :  STD_LOGIC;
                signal tse_pll_s1_grant_vector :  STD_LOGIC;
                signal tse_pll_s1_in_a_read_cycle :  STD_LOGIC;
                signal tse_pll_s1_in_a_write_cycle :  STD_LOGIC;
                signal tse_pll_s1_master_qreq_vector :  STD_LOGIC;
                signal tse_pll_s1_non_bursting_master_requests :  STD_LOGIC;
                signal tse_pll_s1_reg_firsttransfer :  STD_LOGIC;
                signal tse_pll_s1_slavearbiterlockenable :  STD_LOGIC;
                signal tse_pll_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal tse_pll_s1_unreg_firsttransfer :  STD_LOGIC;
                signal tse_pll_s1_waits_for_read :  STD_LOGIC;
                signal tse_pll_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_tse_pll_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT tse_pll_s1_end_xfer;
    end if;

  end process;

  tse_pll_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1);
  --assign tse_pll_s1_readdata_from_sa = tse_pll_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  tse_pll_s1_readdata_from_sa <= tse_pll_s1_readdata;
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1 <= Vector_To_Std_Logic(((std_logic_vector'("00000000000000000000000000000001")) AND (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(((NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read OR NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write)))))));
  --tse_pll_s1_arb_share_counter set values, which is an e_mux
  tse_pll_s1_arb_share_set_values <= std_logic'('1');
  --tse_pll_s1_non_bursting_master_requests mux, which is an e_mux
  tse_pll_s1_non_bursting_master_requests <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1;
  --tse_pll_s1_any_bursting_master_saved_grant mux, which is an e_mux
  tse_pll_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --tse_pll_s1_arb_share_counter_next_value assignment, which is an e_assign
  tse_pll_s1_arb_share_counter_next_value <= Vector_To_Std_Logic(A_WE_StdLogicVector((std_logic'(tse_pll_s1_firsttransfer) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_pll_s1_arb_share_set_values))) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(tse_pll_s1_arb_share_counter) = '1'), (((std_logic_vector'("00000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_pll_s1_arb_share_counter))) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))));
  --tse_pll_s1_allgrants all slave grants, which is an e_mux
  tse_pll_s1_allgrants <= tse_pll_s1_grant_vector;
  --tse_pll_s1_end_xfer assignment, which is an e_assign
  tse_pll_s1_end_xfer <= NOT ((tse_pll_s1_waits_for_read OR tse_pll_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_tse_pll_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_tse_pll_s1 <= tse_pll_s1_end_xfer AND (((NOT tse_pll_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --tse_pll_s1_arb_share_counter arbitration counter enable, which is an e_assign
  tse_pll_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_tse_pll_s1 AND tse_pll_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_tse_pll_s1 AND NOT tse_pll_s1_non_bursting_master_requests));
  --tse_pll_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_pll_s1_arb_share_counter <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'(tse_pll_s1_arb_counter_enable) = '1' then 
        tse_pll_s1_arb_share_counter <= tse_pll_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --tse_pll_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_pll_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((tse_pll_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_tse_pll_s1)) OR ((end_xfer_arb_share_counter_term_tse_pll_s1 AND NOT tse_pll_s1_non_bursting_master_requests)))) = '1' then 
        tse_pll_s1_slavearbiterlockenable <= tse_pll_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/out tse_pll/s1 arbiterlock, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_arbiterlock <= tse_pll_s1_slavearbiterlockenable AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_continuerequest;
  --tse_pll_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  tse_pll_s1_slavearbiterlockenable2 <= tse_pll_s1_arb_share_counter_next_value;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/out tse_pll/s1 arbiterlock2, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_arbiterlock2 <= tse_pll_s1_slavearbiterlockenable2 AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_continuerequest;
  --tse_pll_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  tse_pll_s1_any_continuerequest <= std_logic'('1');
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_continuerequest continued request, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_continuerequest <= std_logic'('1');
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1;
  --tse_pll_s1_writedata mux, which is an e_mux
  tse_pll_s1_writedata <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata;
  --master is always granted when requested
  internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1;
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1/out saved-grant tse_pll/s1, which is an e_assign
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_saved_grant_tse_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1;
  --allow new arb cycle for tse_pll/s1, which is an e_assign
  tse_pll_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  tse_pll_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  tse_pll_s1_master_qreq_vector <= std_logic'('1');
  --tse_pll_s1_reset_n assignment, which is an e_assign
  tse_pll_s1_reset_n <= reset_n;
  --assign tse_pll_s1_resetrequest_from_sa = tse_pll_s1_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  tse_pll_s1_resetrequest_from_sa <= tse_pll_s1_resetrequest;
  tse_pll_s1_chipselect <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1;
  --tse_pll_s1_firsttransfer first transaction, which is an e_assign
  tse_pll_s1_firsttransfer <= A_WE_StdLogic((std_logic'(tse_pll_s1_begins_xfer) = '1'), tse_pll_s1_unreg_firsttransfer, tse_pll_s1_reg_firsttransfer);
  --tse_pll_s1_unreg_firsttransfer first transaction, which is an e_assign
  tse_pll_s1_unreg_firsttransfer <= NOT ((tse_pll_s1_slavearbiterlockenable AND tse_pll_s1_any_continuerequest));
  --tse_pll_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      tse_pll_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(tse_pll_s1_begins_xfer) = '1' then 
        tse_pll_s1_reg_firsttransfer <= tse_pll_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --tse_pll_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  tse_pll_s1_beginbursttransfer_internal <= tse_pll_s1_begins_xfer;
  --tse_pll_s1_read assignment, which is an e_mux
  tse_pll_s1_read <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read;
  --tse_pll_s1_write assignment, which is an e_mux
  tse_pll_s1_write <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write;
  --tse_pll_s1_address mux, which is an e_mux
  tse_pll_s1_address <= NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_nativeaddress;
  --d1_tse_pll_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_tse_pll_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_tse_pll_s1_end_xfer <= tse_pll_s1_end_xfer;
    end if;

  end process;

  --tse_pll_s1_waits_for_read in a cycle, which is an e_mux
  tse_pll_s1_waits_for_read <= tse_pll_s1_in_a_read_cycle AND tse_pll_s1_begins_xfer;
  --tse_pll_s1_in_a_read_cycle assignment, which is an e_assign
  tse_pll_s1_in_a_read_cycle <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read;
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= tse_pll_s1_in_a_read_cycle;
  --tse_pll_s1_waits_for_write in a cycle, which is an e_mux
  tse_pll_s1_waits_for_write <= Vector_To_Std_Logic(((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_pll_s1_in_a_write_cycle))) AND std_logic_vector'("00000000000000000000000000000000")));
  --tse_pll_s1_in_a_write_cycle assignment, which is an e_assign
  tse_pll_s1_in_a_write_cycle <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 AND NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write;
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= tse_pll_s1_in_a_write_cycle;
  wait_for_tse_pll_s1_counter <= std_logic'('0');
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1;
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1;
  --vhdl renameroo for output signals
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1 <= internal_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1;
--synthesis translate_off
    --tse_pll/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity uart1_s1_arbitrator is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                 signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                 signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                 signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal pipeline_bridge_m1_read : IN STD_LOGIC;
                 signal pipeline_bridge_m1_write : IN STD_LOGIC;
                 signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal reset_n : IN STD_LOGIC;
                 signal uart1_s1_dataavailable : IN STD_LOGIC;
                 signal uart1_s1_irq : IN STD_LOGIC;
                 signal uart1_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal uart1_s1_readyfordata : IN STD_LOGIC;

              -- outputs:
                 signal d1_uart1_s1_end_xfer : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_granted_uart1_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_qualified_request_uart1_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_read_data_valid_uart1_s1 : OUT STD_LOGIC;
                 signal pipeline_bridge_m1_requests_uart1_s1 : OUT STD_LOGIC;
                 signal uart1_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                 signal uart1_s1_begintransfer : OUT STD_LOGIC;
                 signal uart1_s1_chipselect : OUT STD_LOGIC;
                 signal uart1_s1_dataavailable_from_sa : OUT STD_LOGIC;
                 signal uart1_s1_irq_from_sa : OUT STD_LOGIC;
                 signal uart1_s1_read_n : OUT STD_LOGIC;
                 signal uart1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal uart1_s1_readyfordata_from_sa : OUT STD_LOGIC;
                 signal uart1_s1_reset_n : OUT STD_LOGIC;
                 signal uart1_s1_write_n : OUT STD_LOGIC;
                 signal uart1_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
              );
end entity uart1_s1_arbitrator;


architecture europa of uart1_s1_arbitrator is
                signal d1_reasons_to_wait :  STD_LOGIC;
                signal enable_nonzero_assertions :  STD_LOGIC;
                signal end_xfer_arb_share_counter_term_uart1_s1 :  STD_LOGIC;
                signal in_a_read_cycle :  STD_LOGIC;
                signal in_a_write_cycle :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_granted_uart1_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_qualified_request_uart1_s1 :  STD_LOGIC;
                signal internal_pipeline_bridge_m1_requests_uart1_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_m1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_m1_continuerequest :  STD_LOGIC;
                signal pipeline_bridge_m1_saved_grant_uart1_s1 :  STD_LOGIC;
                signal shifted_address_to_uart1_s1_from_pipeline_bridge_m1 :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal uart1_s1_allgrants :  STD_LOGIC;
                signal uart1_s1_allow_new_arb_cycle :  STD_LOGIC;
                signal uart1_s1_any_bursting_master_saved_grant :  STD_LOGIC;
                signal uart1_s1_any_continuerequest :  STD_LOGIC;
                signal uart1_s1_arb_counter_enable :  STD_LOGIC;
                signal uart1_s1_arb_share_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal uart1_s1_arb_share_counter_next_value :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal uart1_s1_arb_share_set_values :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal uart1_s1_beginbursttransfer_internal :  STD_LOGIC;
                signal uart1_s1_begins_xfer :  STD_LOGIC;
                signal uart1_s1_end_xfer :  STD_LOGIC;
                signal uart1_s1_firsttransfer :  STD_LOGIC;
                signal uart1_s1_grant_vector :  STD_LOGIC;
                signal uart1_s1_in_a_read_cycle :  STD_LOGIC;
                signal uart1_s1_in_a_write_cycle :  STD_LOGIC;
                signal uart1_s1_master_qreq_vector :  STD_LOGIC;
                signal uart1_s1_non_bursting_master_requests :  STD_LOGIC;
                signal uart1_s1_reg_firsttransfer :  STD_LOGIC;
                signal uart1_s1_slavearbiterlockenable :  STD_LOGIC;
                signal uart1_s1_slavearbiterlockenable2 :  STD_LOGIC;
                signal uart1_s1_unreg_firsttransfer :  STD_LOGIC;
                signal uart1_s1_waits_for_read :  STD_LOGIC;
                signal uart1_s1_waits_for_write :  STD_LOGIC;
                signal wait_for_uart1_s1_counter :  STD_LOGIC;

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_reasons_to_wait <= std_logic'('0');
    elsif clk'event and clk = '1' then
      d1_reasons_to_wait <= NOT uart1_s1_end_xfer;
    end if;

  end process;

  uart1_s1_begins_xfer <= NOT d1_reasons_to_wait AND (internal_pipeline_bridge_m1_qualified_request_uart1_s1);
  --assign uart1_s1_readdata_from_sa = uart1_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart1_s1_readdata_from_sa <= uart1_s1_readdata;
  internal_pipeline_bridge_m1_requests_uart1_s1 <= to_std_logic(((Std_Logic_Vector'(pipeline_bridge_m1_address_to_slave(24 DOWNTO 5) & std_logic_vector'("00000")) = std_logic_vector'("1000000000001100011000000")))) AND pipeline_bridge_m1_chipselect;
  --assign uart1_s1_dataavailable_from_sa = uart1_s1_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart1_s1_dataavailable_from_sa <= uart1_s1_dataavailable;
  --assign uart1_s1_readyfordata_from_sa = uart1_s1_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart1_s1_readyfordata_from_sa <= uart1_s1_readyfordata;
  --uart1_s1_arb_share_counter set values, which is an e_mux
  uart1_s1_arb_share_set_values <= std_logic_vector'("001");
  --uart1_s1_non_bursting_master_requests mux, which is an e_mux
  uart1_s1_non_bursting_master_requests <= internal_pipeline_bridge_m1_requests_uart1_s1;
  --uart1_s1_any_bursting_master_saved_grant mux, which is an e_mux
  uart1_s1_any_bursting_master_saved_grant <= std_logic'('0');
  --uart1_s1_arb_share_counter_next_value assignment, which is an e_assign
  uart1_s1_arb_share_counter_next_value <= A_EXT (A_WE_StdLogicVector((std_logic'(uart1_s1_firsttransfer) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (uart1_s1_arb_share_set_values)) - std_logic_vector'("000000000000000000000000000000001"))), A_WE_StdLogicVector((std_logic'(or_reduce(uart1_s1_arb_share_counter)) = '1'), (((std_logic_vector'("000000000000000000000000000000") & (uart1_s1_arb_share_counter)) - std_logic_vector'("000000000000000000000000000000001"))), std_logic_vector'("000000000000000000000000000000000"))), 3);
  --uart1_s1_allgrants all slave grants, which is an e_mux
  uart1_s1_allgrants <= uart1_s1_grant_vector;
  --uart1_s1_end_xfer assignment, which is an e_assign
  uart1_s1_end_xfer <= NOT ((uart1_s1_waits_for_read OR uart1_s1_waits_for_write));
  --end_xfer_arb_share_counter_term_uart1_s1 arb share counter enable term, which is an e_assign
  end_xfer_arb_share_counter_term_uart1_s1 <= uart1_s1_end_xfer AND (((NOT uart1_s1_any_bursting_master_saved_grant OR in_a_read_cycle) OR in_a_write_cycle));
  --uart1_s1_arb_share_counter arbitration counter enable, which is an e_assign
  uart1_s1_arb_counter_enable <= ((end_xfer_arb_share_counter_term_uart1_s1 AND uart1_s1_allgrants)) OR ((end_xfer_arb_share_counter_term_uart1_s1 AND NOT uart1_s1_non_bursting_master_requests));
  --uart1_s1_arb_share_counter counter, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      uart1_s1_arb_share_counter <= std_logic_vector'("000");
    elsif clk'event and clk = '1' then
      if std_logic'(uart1_s1_arb_counter_enable) = '1' then 
        uart1_s1_arb_share_counter <= uart1_s1_arb_share_counter_next_value;
      end if;
    end if;

  end process;

  --uart1_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      uart1_s1_slavearbiterlockenable <= std_logic'('0');
    elsif clk'event and clk = '1' then
      if std_logic'((((uart1_s1_master_qreq_vector AND end_xfer_arb_share_counter_term_uart1_s1)) OR ((end_xfer_arb_share_counter_term_uart1_s1 AND NOT uart1_s1_non_bursting_master_requests)))) = '1' then 
        uart1_s1_slavearbiterlockenable <= or_reduce(uart1_s1_arb_share_counter_next_value);
      end if;
    end if;

  end process;

  --pipeline_bridge/m1 uart1/s1 arbiterlock, which is an e_assign
  pipeline_bridge_m1_arbiterlock <= uart1_s1_slavearbiterlockenable AND pipeline_bridge_m1_continuerequest;
  --uart1_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  uart1_s1_slavearbiterlockenable2 <= or_reduce(uart1_s1_arb_share_counter_next_value);
  --pipeline_bridge/m1 uart1/s1 arbiterlock2, which is an e_assign
  pipeline_bridge_m1_arbiterlock2 <= uart1_s1_slavearbiterlockenable2 AND pipeline_bridge_m1_continuerequest;
  --uart1_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  uart1_s1_any_continuerequest <= std_logic'('1');
  --pipeline_bridge_m1_continuerequest continued request, which is an e_assign
  pipeline_bridge_m1_continuerequest <= std_logic'('1');
  internal_pipeline_bridge_m1_qualified_request_uart1_s1 <= internal_pipeline_bridge_m1_requests_uart1_s1 AND NOT ((((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect)) AND to_std_logic((((std_logic_vector'("000000000000000000000000000000") & (pipeline_bridge_m1_latency_counter)) /= std_logic_vector'("00000000000000000000000000000000"))))));
  --local readdatavalid pipeline_bridge_m1_read_data_valid_uart1_s1, which is an e_mux
  pipeline_bridge_m1_read_data_valid_uart1_s1 <= (internal_pipeline_bridge_m1_granted_uart1_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))) AND NOT uart1_s1_waits_for_read;
  --uart1_s1_writedata mux, which is an e_mux
  uart1_s1_writedata <= pipeline_bridge_m1_writedata (15 DOWNTO 0);
  --master is always granted when requested
  internal_pipeline_bridge_m1_granted_uart1_s1 <= internal_pipeline_bridge_m1_qualified_request_uart1_s1;
  --pipeline_bridge/m1 saved-grant uart1/s1, which is an e_assign
  pipeline_bridge_m1_saved_grant_uart1_s1 <= internal_pipeline_bridge_m1_requests_uart1_s1;
  --allow new arb cycle for uart1/s1, which is an e_assign
  uart1_s1_allow_new_arb_cycle <= std_logic'('1');
  --placeholder chosen master
  uart1_s1_grant_vector <= std_logic'('1');
  --placeholder vector of master qualified-requests
  uart1_s1_master_qreq_vector <= std_logic'('1');
  uart1_s1_begintransfer <= uart1_s1_begins_xfer;
  --uart1_s1_reset_n assignment, which is an e_assign
  uart1_s1_reset_n <= reset_n;
  uart1_s1_chipselect <= internal_pipeline_bridge_m1_granted_uart1_s1;
  --uart1_s1_firsttransfer first transaction, which is an e_assign
  uart1_s1_firsttransfer <= A_WE_StdLogic((std_logic'(uart1_s1_begins_xfer) = '1'), uart1_s1_unreg_firsttransfer, uart1_s1_reg_firsttransfer);
  --uart1_s1_unreg_firsttransfer first transaction, which is an e_assign
  uart1_s1_unreg_firsttransfer <= NOT ((uart1_s1_slavearbiterlockenable AND uart1_s1_any_continuerequest));
  --uart1_s1_reg_firsttransfer first transaction, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      uart1_s1_reg_firsttransfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      if std_logic'(uart1_s1_begins_xfer) = '1' then 
        uart1_s1_reg_firsttransfer <= uart1_s1_unreg_firsttransfer;
      end if;
    end if;

  end process;

  --uart1_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  uart1_s1_beginbursttransfer_internal <= uart1_s1_begins_xfer;
  --~uart1_s1_read_n assignment, which is an e_mux
  uart1_s1_read_n <= NOT ((internal_pipeline_bridge_m1_granted_uart1_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect))));
  --~uart1_s1_write_n assignment, which is an e_mux
  uart1_s1_write_n <= NOT ((internal_pipeline_bridge_m1_granted_uart1_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect))));
  shifted_address_to_uart1_s1_from_pipeline_bridge_m1 <= pipeline_bridge_m1_address_to_slave;
  --uart1_s1_address mux, which is an e_mux
  uart1_s1_address <= A_EXT (A_SRL(shifted_address_to_uart1_s1_from_pipeline_bridge_m1,std_logic_vector'("00000000000000000000000000000010")), 3);
  --d1_uart1_s1_end_xfer register, which is an e_register
  process (clk, reset_n)
  begin
    if reset_n = '0' then
      d1_uart1_s1_end_xfer <= std_logic'('1');
    elsif clk'event and clk = '1' then
      d1_uart1_s1_end_xfer <= uart1_s1_end_xfer;
    end if;

  end process;

  --uart1_s1_waits_for_read in a cycle, which is an e_mux
  uart1_s1_waits_for_read <= uart1_s1_in_a_read_cycle AND uart1_s1_begins_xfer;
  --uart1_s1_in_a_read_cycle assignment, which is an e_assign
  uart1_s1_in_a_read_cycle <= internal_pipeline_bridge_m1_granted_uart1_s1 AND ((pipeline_bridge_m1_read AND pipeline_bridge_m1_chipselect));
  --in_a_read_cycle assignment, which is an e_mux
  in_a_read_cycle <= uart1_s1_in_a_read_cycle;
  --uart1_s1_waits_for_write in a cycle, which is an e_mux
  uart1_s1_waits_for_write <= uart1_s1_in_a_write_cycle AND uart1_s1_begins_xfer;
  --uart1_s1_in_a_write_cycle assignment, which is an e_assign
  uart1_s1_in_a_write_cycle <= internal_pipeline_bridge_m1_granted_uart1_s1 AND ((pipeline_bridge_m1_write AND pipeline_bridge_m1_chipselect));
  --in_a_write_cycle assignment, which is an e_mux
  in_a_write_cycle <= uart1_s1_in_a_write_cycle;
  wait_for_uart1_s1_counter <= std_logic'('0');
  --assign uart1_s1_irq_from_sa = uart1_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  uart1_s1_irq_from_sa <= uart1_s1_irq;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_granted_uart1_s1 <= internal_pipeline_bridge_m1_granted_uart1_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_qualified_request_uart1_s1 <= internal_pipeline_bridge_m1_qualified_request_uart1_s1;
  --vhdl renameroo for output signals
  pipeline_bridge_m1_requests_uart1_s1 <= internal_pipeline_bridge_m1_requests_uart1_s1;
--synthesis translate_off
    --uart1/s1 enable non-zero assertions, which is an e_register
    process (clk, reset_n)
    begin
      if reset_n = '0' then
        enable_nonzero_assertions <= std_logic'('0');
      elsif clk'event and clk = '1' then
        enable_nonzero_assertions <= std_logic'('1');
      end if;

    end process;

    --pipeline_bridge/m1 non-zero burstcount assertion, which is an e_process
    process (clk)
    VARIABLE write_line64 : line;
    begin
      if clk'event and clk = '1' then
        if std_logic'(((internal_pipeline_bridge_m1_requests_uart1_s1 AND to_std_logic((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pipeline_bridge_m1_burstcount))) = std_logic_vector'("00000000000000000000000000000000"))))) AND enable_nonzero_assertions)) = '1' then 
          write(write_line64, now);
          write(write_line64, string'(": "));
          write(write_line64, string'("pipeline_bridge/m1 drove 0 on its 'burstcount' port while accessing slave uart1/s1"));
          write(output, write_line64.all);
          deallocate (write_line64);
          assert false report "VHDL STOP" severity failure;
        end if;
      end if;

    end process;

--synthesis translate_on

end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_pll_c0_out_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_pll_c0_out_domain_synch_module;


architecture europa of NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_pll_c0_out_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_domain_synch_module;


architecture europa of NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_to_tse_pll_domain_synch_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data_in : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data_out : OUT STD_LOGIC
              );
end entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_to_tse_pll_domain_synch_module;


architecture europa of NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_to_tse_pll_domain_synch_module is
                signal data_in_d1 :  STD_LOGIC;
attribute ALTERA_ATTRIBUTE : string;
attribute ALTERA_ATTRIBUTE of data_in_d1 : signal is "{-from ""*""} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";
attribute ALTERA_ATTRIBUTE of data_out : signal is "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101";

begin

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_in_d1 <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_in_d1 <= data_in;
    end if;

  end process;

  process (clk, reset_n)
  begin
    if reset_n = '0' then
      data_out <= std_logic'('0');
    elsif clk'event and clk = '1' then
      data_out <= data_in_d1;
    end if;

  end process;


end europa;



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc is 
        port (
              -- 1) global signals:
                 signal clk : IN STD_LOGIC;
                 signal clk_to_tse_pll : IN STD_LOGIC;
                 signal pll_c0_out : OUT STD_LOGIC;
                 signal pll_c1_out : OUT STD_LOGIC;
                 signal pll_c2_out : OUT STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal tse_pll_c0_out : OUT STD_LOGIC;

              -- the_button_pio
                 signal in_port_to_the_button_pio : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

              -- the_cpu
                 signal jtag_debug_offchip_trace_clk_from_the_cpu : OUT STD_LOGIC;
                 signal jtag_debug_offchip_trace_data_from_the_cpu : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                 signal jtag_debug_trigout_from_the_cpu : OUT STD_LOGIC;

              -- the_ddr_sdram_0
                 signal clk_to_sdram_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                 signal clk_to_sdram_n_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                 signal ddr_a_from_the_ddr_sdram_0 : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                 signal ddr_ba_from_the_ddr_sdram_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal ddr_cas_n_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                 signal ddr_cke_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                 signal ddr_cs_n_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                 signal ddr_dm_from_the_ddr_sdram_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal ddr_dq_to_and_from_the_ddr_sdram_0 : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                 signal ddr_dqs_to_and_from_the_ddr_sdram_0 : INOUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                 signal ddr_ras_n_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                 signal ddr_we_n_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                 signal dqs_delay_ctrl_to_the_ddr_sdram_0 : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                 signal dqsupdate_to_the_ddr_sdram_0 : IN STD_LOGIC;
                 signal stratix_dll_control_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                 signal write_clk_to_the_ddr_sdram_0 : IN STD_LOGIC;

              -- the_ext_flash_enet_bus_avalon_slave
                 signal ext_flash_enet_bus_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal ext_flash_enet_bus_data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal read_n_to_the_ext_flash : OUT STD_LOGIC;
                 signal select_n_to_the_ext_flash : OUT STD_LOGIC;
                 signal write_n_to_the_ext_flash : OUT STD_LOGIC;

              -- the_ext_ssram_bus_avalon_slave
                 signal adsc_n_to_the_ext_ssram : OUT STD_LOGIC;
                 signal bw_n_to_the_ext_ssram : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal bwe_n_to_the_ext_ssram : OUT STD_LOGIC;
                 signal chipenable1_n_to_the_ext_ssram : OUT STD_LOGIC;
                 signal ext_ssram_bus_address : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                 signal ext_ssram_bus_data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                 signal outputenable_n_to_the_ext_ssram : OUT STD_LOGIC;

              -- the_lcd_display
                 signal LCD_E_from_the_lcd_display : OUT STD_LOGIC;
                 signal LCD_RS_from_the_lcd_display : OUT STD_LOGIC;
                 signal LCD_RW_from_the_lcd_display : OUT STD_LOGIC;
                 signal LCD_data_to_and_from_the_lcd_display : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_led_pio
                 signal out_port_from_the_led_pio : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

              -- the_reconfig_request_pio
                 signal bidir_port_to_and_from_the_reconfig_request_pio : INOUT STD_LOGIC;

              -- the_seven_seg_pio
                 signal out_port_from_the_seven_seg_pio : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

              -- the_tse_mac
                 signal ena_10_from_the_tse_mac : OUT STD_LOGIC;
                 signal eth_mode_from_the_tse_mac : OUT STD_LOGIC;
                 signal gm_rx_d_to_the_tse_mac : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gm_rx_dv_to_the_tse_mac : IN STD_LOGIC;
                 signal gm_rx_err_to_the_tse_mac : IN STD_LOGIC;
                 signal gm_tx_d_from_the_tse_mac : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal gm_tx_en_from_the_tse_mac : OUT STD_LOGIC;
                 signal gm_tx_err_from_the_tse_mac : OUT STD_LOGIC;
                 signal m_rx_col_to_the_tse_mac : IN STD_LOGIC;
                 signal m_rx_crs_to_the_tse_mac : IN STD_LOGIC;
                 signal m_rx_d_to_the_tse_mac : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal m_rx_en_to_the_tse_mac : IN STD_LOGIC;
                 signal m_rx_err_to_the_tse_mac : IN STD_LOGIC;
                 signal m_tx_d_from_the_tse_mac : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal m_tx_en_from_the_tse_mac : OUT STD_LOGIC;
                 signal m_tx_err_from_the_tse_mac : OUT STD_LOGIC;
                 signal mdc_from_the_tse_mac : OUT STD_LOGIC;
                 signal mdio_in_to_the_tse_mac : IN STD_LOGIC;
                 signal mdio_oen_from_the_tse_mac : OUT STD_LOGIC;
                 signal mdio_out_from_the_tse_mac : OUT STD_LOGIC;
                 signal rx_clk_to_the_tse_mac : IN STD_LOGIC;
                 signal set_1000_to_the_tse_mac : IN STD_LOGIC;
                 signal set_10_to_the_tse_mac : IN STD_LOGIC;
                 signal tx_clk_to_the_tse_mac : IN STD_LOGIC;

              -- the_uart1
                 signal rxd_to_the_uart1 : IN STD_LOGIC;
                 signal txd_from_the_uart1 : OUT STD_LOGIC
              );
end entity NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc;


architecture europa of NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc is
component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arbitrator is 
           port (
                 -- inputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_read : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reset_n : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_write : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : OUT STD_LOGIC
                 );
end component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arbitrator;

component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_arbitrator is 
           port (
                 -- inputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_data_valid_pll_s1 : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1 : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_pll_s1_end_xfer : IN STD_LOGIC;
                    signal pll_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_reset_n : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest : OUT STD_LOGIC
                 );
end component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_arbitrator;

component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0;

component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arbitrator is 
           port (
                 -- inputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_read : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reset_n : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_write : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : OUT STD_LOGIC
                 );
end component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arbitrator;

component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_arbitrator is 
           port (
                 -- inputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_data_valid_tse_pll_s1 : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1 : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d1_tse_pll_s1_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal tse_pll_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_reset_n : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest : OUT STD_LOGIC
                 );
end component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_arbitrator;

component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1 is 
           port (
                 -- inputs:
                    signal master_clk : IN STD_LOGIC;
                    signal master_endofpacket : IN STD_LOGIC;
                    signal master_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal master_reset_n : IN STD_LOGIC;
                    signal master_waitrequest : IN STD_LOGIC;
                    signal slave_address : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal slave_byteenable : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal slave_clk : IN STD_LOGIC;
                    signal slave_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal slave_read : IN STD_LOGIC;
                    signal slave_reset_n : IN STD_LOGIC;
                    signal slave_write : IN STD_LOGIC;
                    signal slave_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal master_address : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal master_byteenable : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal master_nativeaddress : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal master_read : OUT STD_LOGIC;
                    signal master_write : OUT STD_LOGIC;
                    signal master_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_endofpacket : OUT STD_LOGIC;
                    signal slave_readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal slave_waitrequest : OUT STD_LOGIC
                 );
end component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1;

component bswap_s1_arbitrator is 
           port (
                 -- inputs:
                    signal bswap_s1_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal bswap_s1_select : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal cpu_custom_instruction_master_combo_dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_custom_instruction_master_combo_datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal bswap_s1_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal bswap_s1_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal bswap_s1_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component bswap_s1_arbitrator;

component bswap is 
           port (
                 -- inputs:
                    signal dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component bswap;

component button_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal button_pio_s1_irq : IN STD_LOGIC;
                    signal button_pio_s1_readdata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal button_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal button_pio_s1_chipselect : OUT STD_LOGIC;
                    signal button_pio_s1_irq_from_sa : OUT STD_LOGIC;
                    signal button_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal button_pio_s1_reset_n : OUT STD_LOGIC;
                    signal button_pio_s1_write_n : OUT STD_LOGIC;
                    signal button_pio_s1_writedata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d1_button_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_button_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_button_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_button_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_button_pio_s1 : OUT STD_LOGIC
                 );
end component button_pio_s1_arbitrator;

component button_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal in_port : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
                 );
end component button_pio;

component cpu_jtag_debug_module_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_jtag_debug_module_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_jtag_debug_module_resetrequest : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_debugaccess : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_jtag_debug_module_address : OUT STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal cpu_jtag_debug_module_begintransfer : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_jtag_debug_module_chipselect : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_debugaccess : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_jtag_debug_module_reset : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_resetrequest_from_sa : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_write : OUT STD_LOGIC;
                    signal cpu_jtag_debug_module_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_cpu_jtag_debug_module_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_cpu_jtag_debug_module : OUT STD_LOGIC
                 );
end component cpu_jtag_debug_module_arbitrator;

component cpu_custom_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal bswap_s1_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal cpu_custom_instruction_master_combo_n : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal interrupt_vector_interrupt_vector_result_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal bswap_s1_select : OUT STD_LOGIC;
                    signal cpu_custom_instruction_master_combo_result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_custom_instruction_master_reset_n : OUT STD_LOGIC;
                    signal interrupt_vector_interrupt_vector_select : OUT STD_LOGIC
                 );
end component cpu_custom_instruction_master_arbitrator;

component cpu_data_master_arbitrator is 
           port (
                 -- inputs:
                    signal button_pio_s1_irq_from_sa : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_granted_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_descriptor_memory_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_ext_ssram_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_packet_memory_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_data_master_granted_tse_mac_control_port : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_ext_ssram_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_packet_memory_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_data_master_qualified_request_tse_mac_control_port : IN STD_LOGIC;
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ext_ssram_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_packet_memory_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_tse_mac_control_port : IN STD_LOGIC;
                    signal cpu_data_master_requests_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_descriptor_memory_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_ext_ssram_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_packet_memory_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_data_master_requests_tse_mac_control_port : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_ddr_sdram_0_s1_end_xfer : IN STD_LOGIC;
                    signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                    signal d1_ext_ssram_bus_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal d1_packet_memory_s1_end_xfer : IN STD_LOGIC;
                    signal d1_pipeline_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal d1_tse_mac_control_port_end_xfer : IN STD_LOGIC;
                    signal ddr_sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ddr_sdram_0_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                    signal descriptor_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal high_res_timer_s1_irq_from_sa : IN STD_LOGIC;
                    signal incoming_ext_ssram_bus_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : IN STD_LOGIC;
                    signal packet_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_csr_irq_from_sa : IN STD_LOGIC;
                    signal sgdma_tx_csr_irq_from_sa : IN STD_LOGIC;
                    signal sys_clk_timer_s1_irq_from_sa : IN STD_LOGIC;
                    signal tse_mac_control_port_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_control_port_waitrequest_from_sa : IN STD_LOGIC;
                    signal uart1_s1_irq_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_data_master_irq : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_data_master_latency_counter : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_data_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_data_master_readdatavalid : OUT STD_LOGIC;
                    signal cpu_data_master_waitrequest : OUT STD_LOGIC
                 );
end component cpu_data_master_arbitrator;

component cpu_instruction_master_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_instruction_master_address : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_instruction_master_granted_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_granted_ext_ssram_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_granted_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_ext_ssram_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_ext_ssram_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_requests_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_requests_ext_ssram_s1 : IN STD_LOGIC;
                    signal cpu_instruction_master_requests_pipeline_bridge_s1 : IN STD_LOGIC;
                    signal d1_ddr_sdram_0_s1_end_xfer : IN STD_LOGIC;
                    signal d1_ext_ssram_bus_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal d1_pipeline_bridge_s1_end_xfer : IN STD_LOGIC;
                    signal ddr_sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ddr_sdram_0_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                    signal incoming_ext_ssram_bus_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_s1_waitrequest_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_instruction_master_address_to_slave : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_instruction_master_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_instruction_master_readdatavalid : OUT STD_LOGIC;
                    signal cpu_instruction_master_waitrequest : OUT STD_LOGIC
                 );
end component cpu_instruction_master_arbitrator;

component cpu is 
           port (
                 -- inputs:
                    signal E_ci_combo_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal d_irq : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d_readdatavalid : IN STD_LOGIC;
                    signal d_waitrequest : IN STD_LOGIC;
                    signal i_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_readdatavalid : IN STD_LOGIC;
                    signal i_waitrequest : IN STD_LOGIC;
                    signal jtag_debug_module_address : IN STD_LOGIC_VECTOR (8 DOWNTO 0);
                    signal jtag_debug_module_begintransfer : IN STD_LOGIC;
                    signal jtag_debug_module_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal jtag_debug_module_clk : IN STD_LOGIC;
                    signal jtag_debug_module_debugaccess : IN STD_LOGIC;
                    signal jtag_debug_module_reset : IN STD_LOGIC;
                    signal jtag_debug_module_select : IN STD_LOGIC;
                    signal jtag_debug_module_write : IN STD_LOGIC;
                    signal jtag_debug_module_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal E_ci_combo_a : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal E_ci_combo_b : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal E_ci_combo_c : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
                    signal E_ci_combo_dataa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal E_ci_combo_datab : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal E_ci_combo_estatus : OUT STD_LOGIC;
                    signal E_ci_combo_ipending : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal E_ci_combo_n : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal E_ci_combo_readra : OUT STD_LOGIC;
                    signal E_ci_combo_readrb : OUT STD_LOGIC;
                    signal E_ci_combo_status : OUT STD_LOGIC;
                    signal E_ci_combo_writerc : OUT STD_LOGIC;
                    signal d_address : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal d_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal d_read : OUT STD_LOGIC;
                    signal d_write : OUT STD_LOGIC;
                    signal d_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal i_address : OUT STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal i_read : OUT STD_LOGIC;
                    signal jtag_debug_module_debugaccess_to_roms : OUT STD_LOGIC;
                    signal jtag_debug_module_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_debug_module_resetrequest : OUT STD_LOGIC;
                    signal jtag_debug_offchip_trace_clk : OUT STD_LOGIC;
                    signal jtag_debug_offchip_trace_data : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal jtag_debug_trigout : OUT STD_LOGIC
                 );
end component cpu;

component ddr_sdram_0_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal ddr_sdram_0_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ddr_sdram_0_s1_readdatavalid : IN STD_LOGIC;
                    signal ddr_sdram_0_s1_waitrequest_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_m_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal sgdma_rx_m_write_write : IN STD_LOGIC;
                    signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal sgdma_tx_m_read_read : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_granted_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_instruction_master_requests_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal d1_ddr_sdram_0_s1_end_xfer : OUT STD_LOGIC;
                    signal ddr_sdram_0_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal ddr_sdram_0_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal ddr_sdram_0_s1_read : OUT STD_LOGIC;
                    signal ddr_sdram_0_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ddr_sdram_0_s1_reset_n : OUT STD_LOGIC;
                    signal ddr_sdram_0_s1_waitrequest_n_from_sa : OUT STD_LOGIC;
                    signal ddr_sdram_0_s1_write : OUT STD_LOGIC;
                    signal ddr_sdram_0_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_m_write_granted_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_m_write_requests_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_granted_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_requests_ddr_sdram_0_s1 : OUT STD_LOGIC
                 );
end component ddr_sdram_0_s1_arbitrator;

component ddr_sdram_0 is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal dqs_delay_ctrl : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal dqsupdate : IN STD_LOGIC;
                    signal local_addr : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal local_be : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal local_read_req : IN STD_LOGIC;
                    signal local_wdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal local_write_req : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_clk : IN STD_LOGIC;

                 -- outputs:
                    signal clk_to_sdram : OUT STD_LOGIC;
                    signal clk_to_sdram_n : OUT STD_LOGIC;
                    signal ddr_a : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal ddr_ba : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ddr_cas_n : OUT STD_LOGIC;
                    signal ddr_cke : OUT STD_LOGIC;
                    signal ddr_cs_n : OUT STD_LOGIC;
                    signal ddr_dm : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ddr_dq : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal ddr_dqs : INOUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ddr_ras_n : OUT STD_LOGIC;
                    signal ddr_we_n : OUT STD_LOGIC;
                    signal local_rdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal local_rdata_valid : OUT STD_LOGIC;
                    signal local_ready : OUT STD_LOGIC;
                    signal stratix_dll_control : OUT STD_LOGIC
                 );
end component ddr_sdram_0;

component descriptor_memory_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_read_latency_counter : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_read : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_write_write : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_read_latency_counter : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_read : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_write_write : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal cpu_data_master_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal d1_descriptor_memory_s1_end_xfer : OUT STD_LOGIC;
                    signal descriptor_memory_s1_address : OUT STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal descriptor_memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal descriptor_memory_s1_chipselect : OUT STD_LOGIC;
                    signal descriptor_memory_s1_clken : OUT STD_LOGIC;
                    signal descriptor_memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_memory_s1_write : OUT STD_LOGIC;
                    signal descriptor_memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_read_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_write_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_write_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_requests_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_write_granted_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_write_requests_descriptor_memory_s1 : OUT STD_LOGIC
                 );
end component descriptor_memory_s1_arbitrator;

component descriptor_memory is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (10 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clken : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component descriptor_memory;

component ext_flash_enet_bus_avalon_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_dbs_address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_dbs_write_8 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_ext_flash_enet_bus_avalon_slave_end_xfer : OUT STD_LOGIC;
                    signal ext_flash_enet_bus_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal ext_flash_enet_bus_data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal ext_flash_s1_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pipeline_bridge_m1_byteenable_ext_flash_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_ext_flash_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_ext_flash_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_ext_flash_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_ext_flash_s1 : OUT STD_LOGIC;
                    signal read_n_to_the_ext_flash : OUT STD_LOGIC;
                    signal select_n_to_the_ext_flash : OUT STD_LOGIC;
                    signal write_n_to_the_ext_flash : OUT STD_LOGIC
                 );
end component ext_flash_enet_bus_avalon_slave_arbitrator;

component ext_flash_enet_bus is 
end component ext_flash_enet_bus;

component ext_flash_enet_bus_bridge_arbitrator is 
end component ext_flash_enet_bus_bridge_arbitrator;

component ext_ssram_bus_avalon_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_m_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal sgdma_rx_m_write_write : IN STD_LOGIC;
                    signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal sgdma_tx_m_read_read : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;

                 -- outputs:
                    signal adsc_n_to_the_ext_ssram : OUT STD_LOGIC;
                    signal bw_n_to_the_ext_ssram : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal bwe_n_to_the_ext_ssram : OUT STD_LOGIC;
                    signal chipenable1_n_to_the_ext_ssram : OUT STD_LOGIC;
                    signal cpu_data_master_granted_ext_ssram_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_ext_ssram_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ext_ssram_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_ext_ssram_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_granted_ext_ssram_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_ext_ssram_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_ext_ssram_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_requests_ext_ssram_s1 : OUT STD_LOGIC;
                    signal d1_ext_ssram_bus_avalon_slave_end_xfer : OUT STD_LOGIC;
                    signal ext_ssram_bus_address : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal ext_ssram_bus_data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal incoming_ext_ssram_bus_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal outputenable_n_to_the_ext_ssram : OUT STD_LOGIC;
                    signal sgdma_rx_m_write_granted_ext_ssram_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_m_write_qualified_request_ext_ssram_s1 : OUT STD_LOGIC;
                    signal sgdma_rx_m_write_requests_ext_ssram_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_granted_ext_ssram_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_qualified_request_ext_ssram_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_ext_ssram_s1 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_requests_ext_ssram_s1 : OUT STD_LOGIC
                 );
end component ext_ssram_bus_avalon_slave_arbitrator;

component ext_ssram_bus is 
end component ext_ssram_bus;

component ext_ssram_bus_bridge_arbitrator is 
end component ext_ssram_bus_bridge_arbitrator;

component high_res_timer_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal high_res_timer_s1_irq : IN STD_LOGIC;
                    signal high_res_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_high_res_timer_s1_end_xfer : OUT STD_LOGIC;
                    signal high_res_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal high_res_timer_s1_chipselect : OUT STD_LOGIC;
                    signal high_res_timer_s1_irq_from_sa : OUT STD_LOGIC;
                    signal high_res_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal high_res_timer_s1_reset_n : OUT STD_LOGIC;
                    signal high_res_timer_s1_write_n : OUT STD_LOGIC;
                    signal high_res_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pipeline_bridge_m1_granted_high_res_timer_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_high_res_timer_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_high_res_timer_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_high_res_timer_s1 : OUT STD_LOGIC
                 );
end component high_res_timer_s1_arbitrator;

component high_res_timer is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component high_res_timer;

component interrupt_vector_interrupt_vector_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_custom_instruction_master_combo_estatus : IN STD_LOGIC;
                    signal cpu_custom_instruction_master_combo_ipending : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal interrupt_vector_interrupt_vector_result : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal interrupt_vector_interrupt_vector_select : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal interrupt_vector_interrupt_vector_estatus : OUT STD_LOGIC;
                    signal interrupt_vector_interrupt_vector_ipending : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal interrupt_vector_interrupt_vector_result_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component interrupt_vector_interrupt_vector_arbitrator;

component interrupt_vector is 
           port (
                 -- inputs:
                    signal estatus : IN STD_LOGIC;
                    signal ipending : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal result : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component interrupt_vector;

component jtag_uart_avalon_jtag_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_dataavailable : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata : IN STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_address : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_chipselect : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_irq_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_read_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_reset_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_write_n : OUT STD_LOGIC;
                    signal jtag_uart_avalon_jtag_slave_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave : OUT STD_LOGIC
                 );
end component jtag_uart_avalon_jtag_slave_arbitrator;

component jtag_uart is 
           port (
                 -- inputs:
                    signal av_address : IN STD_LOGIC;
                    signal av_chipselect : IN STD_LOGIC;
                    signal av_read_n : IN STD_LOGIC;
                    signal av_write_n : IN STD_LOGIC;
                    signal av_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal rst_n : IN STD_LOGIC;

                 -- outputs:
                    signal av_irq : OUT STD_LOGIC;
                    signal av_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal av_waitrequest : OUT STD_LOGIC;
                    signal dataavailable : OUT STD_LOGIC;
                    signal readyfordata : OUT STD_LOGIC
                 );
end component jtag_uart;

component lcd_display_control_slave_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal lcd_display_control_slave_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_lcd_display_control_slave_end_xfer : OUT STD_LOGIC;
                    signal lcd_display_control_slave_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal lcd_display_control_slave_begintransfer : OUT STD_LOGIC;
                    signal lcd_display_control_slave_read : OUT STD_LOGIC;
                    signal lcd_display_control_slave_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal lcd_display_control_slave_wait_counter_eq_0 : OUT STD_LOGIC;
                    signal lcd_display_control_slave_write : OUT STD_LOGIC;
                    signal lcd_display_control_slave_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pipeline_bridge_m1_granted_lcd_display_control_slave : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_lcd_display_control_slave : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_lcd_display_control_slave : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_lcd_display_control_slave : OUT STD_LOGIC
                 );
end component lcd_display_control_slave_arbitrator;

component lcd_display is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal begintransfer : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal LCD_E : OUT STD_LOGIC;
                    signal LCD_RS : OUT STD_LOGIC;
                    signal LCD_RW : OUT STD_LOGIC;
                    signal LCD_data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component lcd_display;

component led_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal led_pio_s1_readdata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_led_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal led_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal led_pio_s1_chipselect : OUT STD_LOGIC;
                    signal led_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal led_pio_s1_reset_n : OUT STD_LOGIC;
                    signal led_pio_s1_write_n : OUT STD_LOGIC;
                    signal led_pio_s1_writedata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pipeline_bridge_m1_granted_led_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_led_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_led_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_led_pio_s1 : OUT STD_LOGIC
                 );
end component led_pio_s1_arbitrator;

component led_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component led_pio;

component packet_memory_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal packet_memory_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_packet_memory_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_packet_memory_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_packet_memory_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_requests_packet_memory_s1 : OUT STD_LOGIC;
                    signal d1_packet_memory_s1_end_xfer : OUT STD_LOGIC;
                    signal packet_memory_s1_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal packet_memory_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal packet_memory_s1_chipselect : OUT STD_LOGIC;
                    signal packet_memory_s1_clken : OUT STD_LOGIC;
                    signal packet_memory_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal packet_memory_s1_write : OUT STD_LOGIC;
                    signal packet_memory_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component packet_memory_s1_arbitrator;

component packet_memory_s2_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal packet_memory_s2_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_m_write_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal sgdma_rx_m_write_write : IN STD_LOGIC;
                    signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_address_to_slave : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal sgdma_tx_m_read_read : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;

                 -- outputs:
                    signal d1_packet_memory_s2_end_xfer : OUT STD_LOGIC;
                    signal packet_memory_s2_address : OUT STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal packet_memory_s2_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal packet_memory_s2_chipselect : OUT STD_LOGIC;
                    signal packet_memory_s2_clken : OUT STD_LOGIC;
                    signal packet_memory_s2_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal packet_memory_s2_write : OUT STD_LOGIC;
                    signal packet_memory_s2_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_m_write_granted_packet_memory_s2 : OUT STD_LOGIC;
                    signal sgdma_rx_m_write_qualified_request_packet_memory_s2 : OUT STD_LOGIC;
                    signal sgdma_rx_m_write_requests_packet_memory_s2 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_granted_packet_memory_s2 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_qualified_request_packet_memory_s2 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_packet_memory_s2 : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_requests_packet_memory_s2 : OUT STD_LOGIC
                 );
end component packet_memory_s2_arbitrator;

component packet_memory is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal address2 : IN STD_LOGIC_VECTOR (13 DOWNTO 0);
                    signal byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal byteenable2 : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal chipselect2 : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal clk2 : IN STD_LOGIC;
                    signal clken : IN STD_LOGIC;
                    signal clken2 : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal write2 : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal writedata2 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal readdata2 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component packet_memory;

component pipeline_bridge_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_data_master_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal cpu_data_master_debugaccess : IN STD_LOGIC;
                    signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal cpu_instruction_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_instruction_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_instruction_master_read : IN STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal pipeline_bridge_s1_endofpacket : IN STD_LOGIC;
                    signal pipeline_bridge_s1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_s1_readdatavalid : IN STD_LOGIC;
                    signal pipeline_bridge_s1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_data_master_requests_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_granted_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_qualified_request_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register : OUT STD_LOGIC;
                    signal cpu_instruction_master_requests_pipeline_bridge_s1 : OUT STD_LOGIC;
                    signal d1_pipeline_bridge_s1_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_address : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal pipeline_bridge_s1_arbiterlock : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_arbiterlock2 : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_burstcount : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_s1_chipselect : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_debugaccess : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_endofpacket_from_sa : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_nativeaddress : OUT STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal pipeline_bridge_s1_read : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_s1_reset_n : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_waitrequest_from_sa : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_write : OUT STD_LOGIC;
                    signal pipeline_bridge_s1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component pipeline_bridge_s1_arbitrator;

component pipeline_bridge_m1_arbitrator is 
           port (
                 -- inputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa : IN STD_LOGIC;
                    signal button_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal cpu_jtag_debug_module_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer : IN STD_LOGIC;
                    signal d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer : IN STD_LOGIC;
                    signal d1_button_pio_s1_end_xfer : IN STD_LOGIC;
                    signal d1_cpu_jtag_debug_module_end_xfer : IN STD_LOGIC;
                    signal d1_ext_flash_enet_bus_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal d1_high_res_timer_s1_end_xfer : IN STD_LOGIC;
                    signal d1_jtag_uart_avalon_jtag_slave_end_xfer : IN STD_LOGIC;
                    signal d1_lcd_display_control_slave_end_xfer : IN STD_LOGIC;
                    signal d1_led_pio_s1_end_xfer : IN STD_LOGIC;
                    signal d1_reconfig_request_pio_s1_end_xfer : IN STD_LOGIC;
                    signal d1_seven_seg_pio_s1_end_xfer : IN STD_LOGIC;
                    signal d1_sgdma_rx_csr_end_xfer : IN STD_LOGIC;
                    signal d1_sgdma_tx_csr_end_xfer : IN STD_LOGIC;
                    signal d1_sys_clk_timer_s1_end_xfer : IN STD_LOGIC;
                    signal d1_uart1_s1_end_xfer : IN STD_LOGIC;
                    signal ext_flash_s1_wait_counter_eq_0 : IN STD_LOGIC;
                    signal high_res_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa : IN STD_LOGIC;
                    signal lcd_display_control_slave_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal lcd_display_control_slave_wait_counter_eq_0 : IN STD_LOGIC;
                    signal led_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pipeline_bridge_m1_address : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal pipeline_bridge_m1_byteenable_ext_flash_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_button_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_ext_flash_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_high_res_timer_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_lcd_display_control_slave : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_led_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_reconfig_request_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_seven_seg_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_sgdma_rx_csr : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_sgdma_tx_csr : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_granted_uart1_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_button_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_ext_flash_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_high_res_timer_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_lcd_display_control_slave : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_led_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_sgdma_rx_csr : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_sgdma_tx_csr : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_uart1_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_button_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_ext_flash_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_high_res_timer_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_lcd_display_control_slave : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_led_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_sgdma_rx_csr : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_sgdma_tx_csr : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_uart1_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_button_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_cpu_jtag_debug_module : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_ext_flash_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_high_res_timer_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_lcd_display_control_slave : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_led_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_reconfig_request_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_seven_seg_pio_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_sgdma_rx_csr : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_sgdma_tx_csr : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_sys_clk_timer_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_requests_uart1_s1 : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reconfig_request_pio_s1_readdata_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal seven_seg_pio_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sgdma_rx_csr_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_csr_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sys_clk_timer_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal uart1_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal pipeline_bridge_m1_address_to_slave : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_dbs_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_dbs_write_8 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal pipeline_bridge_m1_endofpacket : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal pipeline_bridge_m1_readdatavalid : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_waitrequest : OUT STD_LOGIC
                 );
end component pipeline_bridge_m1_arbitrator;

component pipeline_bridge is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal m1_endofpacket : IN STD_LOGIC;
                    signal m1_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m1_readdatavalid : IN STD_LOGIC;
                    signal m1_waitrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal s1_address : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal s1_arbiterlock : IN STD_LOGIC;
                    signal s1_arbiterlock2 : IN STD_LOGIC;
                    signal s1_burstcount : IN STD_LOGIC;
                    signal s1_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal s1_chipselect : IN STD_LOGIC;
                    signal s1_debugaccess : IN STD_LOGIC;
                    signal s1_nativeaddress : IN STD_LOGIC_VECTOR (22 DOWNTO 0);
                    signal s1_read : IN STD_LOGIC;
                    signal s1_write : IN STD_LOGIC;
                    signal s1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal m1_address : OUT STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal m1_burstcount : OUT STD_LOGIC;
                    signal m1_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m1_chipselect : OUT STD_LOGIC;
                    signal m1_debugaccess : OUT STD_LOGIC;
                    signal m1_read : OUT STD_LOGIC;
                    signal m1_write : OUT STD_LOGIC;
                    signal m1_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal s1_endofpacket : OUT STD_LOGIC;
                    signal s1_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal s1_readdatavalid : OUT STD_LOGIC;
                    signal s1_waitrequest : OUT STD_LOGIC
                 );
end component pipeline_bridge;

component pipeline_bridge_bridge_arbitrator is 
end component pipeline_bridge_bridge_arbitrator;

component pll_s1_arbitrator is 
           port (
                 -- inputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal pll_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pll_s1_resetrequest : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_data_valid_pll_s1 : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1 : OUT STD_LOGIC;
                    signal d1_pll_s1_end_xfer : OUT STD_LOGIC;
                    signal pll_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal pll_s1_chipselect : OUT STD_LOGIC;
                    signal pll_s1_read : OUT STD_LOGIC;
                    signal pll_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal pll_s1_reset_n : OUT STD_LOGIC;
                    signal pll_s1_resetrequest_from_sa : OUT STD_LOGIC;
                    signal pll_s1_write : OUT STD_LOGIC;
                    signal pll_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component pll_s1_arbitrator;

component pll is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal c0 : OUT STD_LOGIC;
                    signal c1 : OUT STD_LOGIC;
                    signal c2 : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal resetrequest : OUT STD_LOGIC
                 );
end component pll;

component reconfig_request_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reconfig_request_pio_s1_readdata : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal d1_reconfig_request_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_reconfig_request_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_reconfig_request_pio_s1 : OUT STD_LOGIC;
                    signal reconfig_request_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal reconfig_request_pio_s1_chipselect : OUT STD_LOGIC;
                    signal reconfig_request_pio_s1_readdata_from_sa : OUT STD_LOGIC;
                    signal reconfig_request_pio_s1_reset_n : OUT STD_LOGIC;
                    signal reconfig_request_pio_s1_write_n : OUT STD_LOGIC;
                    signal reconfig_request_pio_s1_writedata : OUT STD_LOGIC
                 );
end component reconfig_request_pio_s1_arbitrator;

component reconfig_request_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC;

                 -- outputs:
                    signal bidir_port : INOUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC
                 );
end component reconfig_request_pio;

component seven_seg_pio_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal seven_seg_pio_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal d1_seven_seg_pio_s1_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_seven_seg_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_seven_seg_pio_s1 : OUT STD_LOGIC;
                    signal seven_seg_pio_s1_address : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal seven_seg_pio_s1_chipselect : OUT STD_LOGIC;
                    signal seven_seg_pio_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal seven_seg_pio_s1_reset_n : OUT STD_LOGIC;
                    signal seven_seg_pio_s1_write_n : OUT STD_LOGIC;
                    signal seven_seg_pio_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component seven_seg_pio_s1_arbitrator;

component seven_seg_pio is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal out_port : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component seven_seg_pio;

component sgdma_rx_csr_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_csr_irq : IN STD_LOGIC;
                    signal sgdma_rx_csr_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal d1_sgdma_rx_csr_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_sgdma_rx_csr : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_sgdma_rx_csr : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_sgdma_rx_csr : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_sgdma_rx_csr : OUT STD_LOGIC;
                    signal sgdma_rx_csr_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal sgdma_rx_csr_chipselect : OUT STD_LOGIC;
                    signal sgdma_rx_csr_irq_from_sa : OUT STD_LOGIC;
                    signal sgdma_rx_csr_read : OUT STD_LOGIC;
                    signal sgdma_rx_csr_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_csr_reset_n : OUT STD_LOGIC;
                    signal sgdma_rx_csr_write : OUT STD_LOGIC;
                    signal sgdma_rx_csr_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sgdma_rx_csr_arbitrator;

component sgdma_rx_in_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_in_ready : IN STD_LOGIC;
                    signal tse_mac_receive_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_receive_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal tse_mac_receive_endofpacket : IN STD_LOGIC;
                    signal tse_mac_receive_error : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal tse_mac_receive_startofpacket : IN STD_LOGIC;
                    signal tse_mac_receive_valid : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_rx_in_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_in_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sgdma_rx_in_endofpacket : OUT STD_LOGIC;
                    signal sgdma_rx_in_error : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal sgdma_rx_in_ready_from_sa : OUT STD_LOGIC;
                    signal sgdma_rx_in_startofpacket : OUT STD_LOGIC;
                    signal sgdma_rx_in_valid : OUT STD_LOGIC
                 );
end component sgdma_rx_in_arbitrator;

component sgdma_rx_descriptor_read_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                    signal descriptor_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_read_granted_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_read : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_read_requests_descriptor_memory_s1 : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_rx_descriptor_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_read_latency_counter : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_read_readdatavalid : OUT STD_LOGIC;
                    signal sgdma_rx_descriptor_read_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_rx_descriptor_read_arbitrator;

component sgdma_rx_descriptor_write_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_write_granted_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_requests_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_write : IN STD_LOGIC;
                    signal sgdma_rx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal sgdma_rx_descriptor_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_descriptor_write_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_rx_descriptor_write_arbitrator;

component sgdma_rx_m_write_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_ddr_sdram_0_s1_end_xfer : IN STD_LOGIC;
                    signal d1_ext_ssram_bus_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal d1_packet_memory_s2_end_xfer : IN STD_LOGIC;
                    signal ddr_sdram_0_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_m_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_m_write_byteenable : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal sgdma_rx_m_write_granted_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_granted_ext_ssram_s1 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_granted_packet_memory_s2 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_qualified_request_ext_ssram_s1 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_qualified_request_packet_memory_s2 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_requests_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_requests_ext_ssram_s1 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_requests_packet_memory_s2 : IN STD_LOGIC;
                    signal sgdma_rx_m_write_write : IN STD_LOGIC;
                    signal sgdma_rx_m_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal sgdma_rx_m_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_rx_m_write_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_rx_m_write_arbitrator;

component sgdma_rx is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal csr_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal csr_chipselect : IN STD_LOGIC;
                    signal csr_read : IN STD_LOGIC;
                    signal csr_write : IN STD_LOGIC;
                    signal csr_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_readdatavalid : IN STD_LOGIC;
                    signal descriptor_read_waitrequest : IN STD_LOGIC;
                    signal descriptor_write_waitrequest : IN STD_LOGIC;
                    signal in_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal in_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal in_endofpacket : IN STD_LOGIC;
                    signal in_error : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal in_startofpacket : IN STD_LOGIC;
                    signal in_valid : IN STD_LOGIC;
                    signal m_write_waitrequest : IN STD_LOGIC;
                    signal system_reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal csr_irq : OUT STD_LOGIC;
                    signal csr_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_read : OUT STD_LOGIC;
                    signal descriptor_write_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_write_write : OUT STD_LOGIC;
                    signal descriptor_write_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal in_ready : OUT STD_LOGIC;
                    signal m_write_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m_write_byteenable : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_write_write : OUT STD_LOGIC;
                    signal m_write_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sgdma_rx;

component sgdma_tx_csr_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_csr_irq : IN STD_LOGIC;
                    signal sgdma_tx_csr_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal d1_sgdma_tx_csr_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_sgdma_tx_csr : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_sgdma_tx_csr : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_sgdma_tx_csr : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_sgdma_tx_csr : OUT STD_LOGIC;
                    signal sgdma_tx_csr_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal sgdma_tx_csr_chipselect : OUT STD_LOGIC;
                    signal sgdma_tx_csr_irq_from_sa : OUT STD_LOGIC;
                    signal sgdma_tx_csr_read : OUT STD_LOGIC;
                    signal sgdma_tx_csr_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_csr_reset_n : OUT STD_LOGIC;
                    signal sgdma_tx_csr_write : OUT STD_LOGIC;
                    signal sgdma_tx_csr_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component sgdma_tx_csr_arbitrator;

component sgdma_tx_descriptor_read_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                    signal descriptor_memory_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_read_granted_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_read : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_read_requests_descriptor_memory_s1 : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_tx_descriptor_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_read_latency_counter : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_read_readdatavalid : OUT STD_LOGIC;
                    signal sgdma_tx_descriptor_read_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_tx_descriptor_read_arbitrator;

component sgdma_tx_descriptor_write_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_descriptor_memory_s1_end_xfer : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_write_granted_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_requests_descriptor_memory_s1 : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_write : IN STD_LOGIC;
                    signal sgdma_tx_descriptor_write_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal sgdma_tx_descriptor_write_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_descriptor_write_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_tx_descriptor_write_arbitrator;

component sgdma_tx_m_read_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal d1_ddr_sdram_0_s1_end_xfer : IN STD_LOGIC;
                    signal d1_ext_ssram_bus_avalon_slave_end_xfer : IN STD_LOGIC;
                    signal d1_packet_memory_s2_end_xfer : IN STD_LOGIC;
                    signal ddr_sdram_0_s1_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ddr_sdram_0_s1_waitrequest_n_from_sa : IN STD_LOGIC;
                    signal incoming_ext_ssram_bus_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal packet_memory_s2_readdata_from_sa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_m_read_address : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_granted_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_granted_ext_ssram_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_granted_packet_memory_s2 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_qualified_request_ext_ssram_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_qualified_request_packet_memory_s2 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_ext_ssram_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_read_data_valid_packet_memory_s2 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_requests_ddr_sdram_0_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_requests_ext_ssram_s1 : IN STD_LOGIC;
                    signal sgdma_tx_m_read_requests_packet_memory_s2 : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_tx_m_read_address_to_slave : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_latency_counter : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal sgdma_tx_m_read_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_m_read_readdatavalid : OUT STD_LOGIC;
                    signal sgdma_tx_m_read_waitrequest : OUT STD_LOGIC
                 );
end component sgdma_tx_m_read_arbitrator;

component sgdma_tx_out_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sgdma_tx_out_endofpacket : IN STD_LOGIC;
                    signal sgdma_tx_out_error : IN STD_LOGIC;
                    signal sgdma_tx_out_startofpacket : IN STD_LOGIC;
                    signal sgdma_tx_out_valid : IN STD_LOGIC;
                    signal tse_mac_transmit_ready_from_sa : IN STD_LOGIC;

                 -- outputs:
                    signal sgdma_tx_out_ready : OUT STD_LOGIC
                 );
end component sgdma_tx_out_arbitrator;

component sgdma_tx is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal csr_address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal csr_chipselect : IN STD_LOGIC;
                    signal csr_read : IN STD_LOGIC;
                    signal csr_write : IN STD_LOGIC;
                    signal csr_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_readdatavalid : IN STD_LOGIC;
                    signal descriptor_read_waitrequest : IN STD_LOGIC;
                    signal descriptor_write_waitrequest : IN STD_LOGIC;
                    signal m_read_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m_read_readdatavalid : IN STD_LOGIC;
                    signal m_read_waitrequest : IN STD_LOGIC;
                    signal out_ready : IN STD_LOGIC;
                    signal system_reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal csr_irq : OUT STD_LOGIC;
                    signal csr_readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_read_read : OUT STD_LOGIC;
                    signal descriptor_write_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal descriptor_write_write : OUT STD_LOGIC;
                    signal descriptor_write_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m_read_address : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal m_read_read : OUT STD_LOGIC;
                    signal out_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal out_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal out_endofpacket : OUT STD_LOGIC;
                    signal out_error : OUT STD_LOGIC;
                    signal out_startofpacket : OUT STD_LOGIC;
                    signal out_valid : OUT STD_LOGIC
                 );
end component sgdma_tx;

component sys_clk_timer_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal sys_clk_timer_s1_irq : IN STD_LOGIC;
                    signal sys_clk_timer_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal d1_sys_clk_timer_s1_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_sys_clk_timer_s1 : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal sys_clk_timer_s1_chipselect : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_irq_from_sa : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal sys_clk_timer_s1_reset_n : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_write_n : OUT STD_LOGIC;
                    signal sys_clk_timer_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sys_clk_timer_s1_arbitrator;

component sys_clk_timer is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component sys_clk_timer;

component tse_mac_control_port_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal cpu_data_master_address_to_slave : IN STD_LOGIC_VECTOR (27 DOWNTO 0);
                    signal cpu_data_master_latency_counter : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal cpu_data_master_read : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register : IN STD_LOGIC;
                    signal cpu_data_master_write : IN STD_LOGIC;
                    signal cpu_data_master_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal tse_mac_control_port_readdata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_control_port_waitrequest : IN STD_LOGIC;

                 -- outputs:
                    signal cpu_data_master_granted_tse_mac_control_port : OUT STD_LOGIC;
                    signal cpu_data_master_qualified_request_tse_mac_control_port : OUT STD_LOGIC;
                    signal cpu_data_master_read_data_valid_tse_mac_control_port : OUT STD_LOGIC;
                    signal cpu_data_master_requests_tse_mac_control_port : OUT STD_LOGIC;
                    signal d1_tse_mac_control_port_end_xfer : OUT STD_LOGIC;
                    signal tse_mac_control_port_address : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal tse_mac_control_port_read : OUT STD_LOGIC;
                    signal tse_mac_control_port_readdata_from_sa : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_control_port_reset : OUT STD_LOGIC;
                    signal tse_mac_control_port_waitrequest_from_sa : OUT STD_LOGIC;
                    signal tse_mac_control_port_write : OUT STD_LOGIC;
                    signal tse_mac_control_port_writedata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component tse_mac_control_port_arbitrator;

component tse_mac_transmit_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_tx_out_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal sgdma_tx_out_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal sgdma_tx_out_endofpacket : IN STD_LOGIC;
                    signal sgdma_tx_out_error : IN STD_LOGIC;
                    signal sgdma_tx_out_startofpacket : IN STD_LOGIC;
                    signal sgdma_tx_out_valid : IN STD_LOGIC;
                    signal tse_mac_transmit_ready : IN STD_LOGIC;

                 -- outputs:
                    signal tse_mac_transmit_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_transmit_empty : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal tse_mac_transmit_endofpacket : OUT STD_LOGIC;
                    signal tse_mac_transmit_error : OUT STD_LOGIC;
                    signal tse_mac_transmit_ready_from_sa : OUT STD_LOGIC;
                    signal tse_mac_transmit_startofpacket : OUT STD_LOGIC;
                    signal tse_mac_transmit_valid : OUT STD_LOGIC
                 );
end component tse_mac_transmit_arbitrator;

component tse_mac_receive_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal sgdma_rx_in_ready_from_sa : IN STD_LOGIC;
                    signal tse_mac_receive_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal tse_mac_receive_empty : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal tse_mac_receive_endofpacket : IN STD_LOGIC;
                    signal tse_mac_receive_error : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal tse_mac_receive_startofpacket : IN STD_LOGIC;
                    signal tse_mac_receive_valid : IN STD_LOGIC;

                 -- outputs:
                    signal tse_mac_receive_ready : OUT STD_LOGIC
                 );
end component tse_mac_receive_arbitrator;

component tse_mac is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal ff_rx_clk : IN STD_LOGIC;
                    signal ff_rx_rdy : IN STD_LOGIC;
                    signal ff_tx_clk : IN STD_LOGIC;
                    signal ff_tx_data : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ff_tx_eop : IN STD_LOGIC;
                    signal ff_tx_err : IN STD_LOGIC;
                    signal ff_tx_mod : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ff_tx_sop : IN STD_LOGIC;
                    signal ff_tx_wren : IN STD_LOGIC;
                    signal gm_rx_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_rx_dv : IN STD_LOGIC;
                    signal gm_rx_err : IN STD_LOGIC;
                    signal m_rx_col : IN STD_LOGIC;
                    signal m_rx_crs : IN STD_LOGIC;
                    signal m_rx_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_rx_en : IN STD_LOGIC;
                    signal m_rx_err : IN STD_LOGIC;
                    signal mdio_in : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset : IN STD_LOGIC;
                    signal rx_clk : IN STD_LOGIC;
                    signal set_10 : IN STD_LOGIC;
                    signal set_1000 : IN STD_LOGIC;
                    signal tx_clk : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);

                 -- outputs:
                    signal ena_10 : OUT STD_LOGIC;
                    signal eth_mode : OUT STD_LOGIC;
                    signal ff_rx_data : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal ff_rx_dval : OUT STD_LOGIC;
                    signal ff_rx_eop : OUT STD_LOGIC;
                    signal ff_rx_mod : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ff_rx_sop : OUT STD_LOGIC;
                    signal ff_tx_rdy : OUT STD_LOGIC;
                    signal gm_tx_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_tx_en : OUT STD_LOGIC;
                    signal gm_tx_err : OUT STD_LOGIC;
                    signal m_tx_d : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_tx_en : OUT STD_LOGIC;
                    signal m_tx_err : OUT STD_LOGIC;
                    signal mdc : OUT STD_LOGIC;
                    signal mdio_oen : OUT STD_LOGIC;
                    signal mdio_out : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal rx_err : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal waitrequest : OUT STD_LOGIC
                 );
end component tse_mac;

component tse_pll_s1_arbitrator is 
           port (
                 -- inputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_nativeaddress : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write : IN STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal clk : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal tse_pll_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal tse_pll_s1_resetrequest : IN STD_LOGIC;

                 -- outputs:
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_data_valid_tse_pll_s1 : OUT STD_LOGIC;
                    signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1 : OUT STD_LOGIC;
                    signal d1_tse_pll_s1_end_xfer : OUT STD_LOGIC;
                    signal tse_pll_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal tse_pll_s1_chipselect : OUT STD_LOGIC;
                    signal tse_pll_s1_read : OUT STD_LOGIC;
                    signal tse_pll_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal tse_pll_s1_reset_n : OUT STD_LOGIC;
                    signal tse_pll_s1_resetrequest_from_sa : OUT STD_LOGIC;
                    signal tse_pll_s1_write : OUT STD_LOGIC;
                    signal tse_pll_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component tse_pll_s1_arbitrator;

component tse_pll is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal write : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal c0 : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal resetrequest : OUT STD_LOGIC
                 );
end component tse_pll;

component uart1_s1_arbitrator is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal pipeline_bridge_m1_address_to_slave : IN STD_LOGIC_VECTOR (24 DOWNTO 0);
                    signal pipeline_bridge_m1_burstcount : IN STD_LOGIC;
                    signal pipeline_bridge_m1_chipselect : IN STD_LOGIC;
                    signal pipeline_bridge_m1_latency_counter : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal pipeline_bridge_m1_read : IN STD_LOGIC;
                    signal pipeline_bridge_m1_write : IN STD_LOGIC;
                    signal pipeline_bridge_m1_writedata : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal reset_n : IN STD_LOGIC;
                    signal uart1_s1_dataavailable : IN STD_LOGIC;
                    signal uart1_s1_irq : IN STD_LOGIC;
                    signal uart1_s1_readdata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal uart1_s1_readyfordata : IN STD_LOGIC;

                 -- outputs:
                    signal d1_uart1_s1_end_xfer : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_granted_uart1_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_qualified_request_uart1_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_read_data_valid_uart1_s1 : OUT STD_LOGIC;
                    signal pipeline_bridge_m1_requests_uart1_s1 : OUT STD_LOGIC;
                    signal uart1_s1_address : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal uart1_s1_begintransfer : OUT STD_LOGIC;
                    signal uart1_s1_chipselect : OUT STD_LOGIC;
                    signal uart1_s1_dataavailable_from_sa : OUT STD_LOGIC;
                    signal uart1_s1_irq_from_sa : OUT STD_LOGIC;
                    signal uart1_s1_read_n : OUT STD_LOGIC;
                    signal uart1_s1_readdata_from_sa : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal uart1_s1_readyfordata_from_sa : OUT STD_LOGIC;
                    signal uart1_s1_reset_n : OUT STD_LOGIC;
                    signal uart1_s1_write_n : OUT STD_LOGIC;
                    signal uart1_s1_writedata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
                 );
end component uart1_s1_arbitrator;

component uart1 is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
                    signal begintransfer : IN STD_LOGIC;
                    signal chipselect : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal read_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal rxd : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;
                    signal writedata : IN STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- outputs:
                    signal dataavailable : OUT STD_LOGIC;
                    signal irq : OUT STD_LOGIC;
                    signal readdata : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal readyfordata : OUT STD_LOGIC;
                    signal txd : OUT STD_LOGIC
                 );
end component uart1;

component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_pll_c0_out_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_pll_c0_out_domain_synch_module;

component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_domain_synch_module;

component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_to_tse_pll_domain_synch_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data_in : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data_out : OUT STD_LOGIC
                 );
end component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_to_tse_pll_domain_synch_module;

                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_read :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reset_n :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_write :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_endofpacket :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_data_valid_pll_s1 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_reset_n :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_read :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reset_n :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_write :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_endofpacket :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_nativeaddress :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_data_valid_tse_pll_s1 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1 :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_reset_n :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal bswap_s1_dataa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal bswap_s1_datab :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal bswap_s1_result :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal bswap_s1_result_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal bswap_s1_select :  STD_LOGIC;
                signal button_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal button_pio_s1_chipselect :  STD_LOGIC;
                signal button_pio_s1_irq :  STD_LOGIC;
                signal button_pio_s1_irq_from_sa :  STD_LOGIC;
                signal button_pio_s1_readdata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal button_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal button_pio_s1_reset_n :  STD_LOGIC;
                signal button_pio_s1_write_n :  STD_LOGIC;
                signal button_pio_s1_writedata :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal clk_reset_n :  STD_LOGIC;
                signal clk_to_tse_pll_reset_n :  STD_LOGIC;
                signal cpu_custom_instruction_master_combo_a :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_b :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_c :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_dataa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_datab :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_estatus :  STD_LOGIC;
                signal cpu_custom_instruction_master_combo_ipending :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_n :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_readra :  STD_LOGIC;
                signal cpu_custom_instruction_master_combo_readrb :  STD_LOGIC;
                signal cpu_custom_instruction_master_combo_result :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_status :  STD_LOGIC;
                signal cpu_custom_instruction_master_combo_writerc :  STD_LOGIC;
                signal cpu_custom_instruction_master_reset_n :  STD_LOGIC;
                signal cpu_data_master_address :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_data_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_data_master_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_data_master_debugaccess :  STD_LOGIC;
                signal cpu_data_master_granted_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_ext_ssram_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_packet_memory_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_data_master_granted_tse_mac_control_port :  STD_LOGIC;
                signal cpu_data_master_irq :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_data_master_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal cpu_data_master_qualified_request_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_ext_ssram_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_packet_memory_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_data_master_qualified_request_tse_mac_control_port :  STD_LOGIC;
                signal cpu_data_master_read :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_descriptor_memory_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_ext_ssram_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_packet_memory_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register :  STD_LOGIC;
                signal cpu_data_master_read_data_valid_tse_mac_control_port :  STD_LOGIC;
                signal cpu_data_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_data_master_readdatavalid :  STD_LOGIC;
                signal cpu_data_master_requests_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_ext_ssram_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_packet_memory_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_data_master_requests_tse_mac_control_port :  STD_LOGIC;
                signal cpu_data_master_waitrequest :  STD_LOGIC;
                signal cpu_data_master_write :  STD_LOGIC;
                signal cpu_data_master_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_instruction_master_address :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_instruction_master_address_to_slave :  STD_LOGIC_VECTOR (27 DOWNTO 0);
                signal cpu_instruction_master_granted_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_instruction_master_granted_ext_ssram_s1 :  STD_LOGIC;
                signal cpu_instruction_master_granted_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_instruction_master_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal cpu_instruction_master_qualified_request_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_instruction_master_qualified_request_ext_ssram_s1 :  STD_LOGIC;
                signal cpu_instruction_master_qualified_request_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_instruction_master_read :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_ext_ssram_s1 :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register :  STD_LOGIC;
                signal cpu_instruction_master_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_instruction_master_readdatavalid :  STD_LOGIC;
                signal cpu_instruction_master_requests_ddr_sdram_0_s1 :  STD_LOGIC;
                signal cpu_instruction_master_requests_ext_ssram_s1 :  STD_LOGIC;
                signal cpu_instruction_master_requests_pipeline_bridge_s1 :  STD_LOGIC;
                signal cpu_instruction_master_waitrequest :  STD_LOGIC;
                signal cpu_jtag_debug_module_address :  STD_LOGIC_VECTOR (8 DOWNTO 0);
                signal cpu_jtag_debug_module_begintransfer :  STD_LOGIC;
                signal cpu_jtag_debug_module_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal cpu_jtag_debug_module_chipselect :  STD_LOGIC;
                signal cpu_jtag_debug_module_debugaccess :  STD_LOGIC;
                signal cpu_jtag_debug_module_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_jtag_debug_module_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal cpu_jtag_debug_module_reset :  STD_LOGIC;
                signal cpu_jtag_debug_module_resetrequest :  STD_LOGIC;
                signal cpu_jtag_debug_module_resetrequest_from_sa :  STD_LOGIC;
                signal cpu_jtag_debug_module_write :  STD_LOGIC;
                signal cpu_jtag_debug_module_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer :  STD_LOGIC;
                signal d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer :  STD_LOGIC;
                signal d1_button_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_cpu_jtag_debug_module_end_xfer :  STD_LOGIC;
                signal d1_ddr_sdram_0_s1_end_xfer :  STD_LOGIC;
                signal d1_descriptor_memory_s1_end_xfer :  STD_LOGIC;
                signal d1_ext_flash_enet_bus_avalon_slave_end_xfer :  STD_LOGIC;
                signal d1_ext_ssram_bus_avalon_slave_end_xfer :  STD_LOGIC;
                signal d1_high_res_timer_s1_end_xfer :  STD_LOGIC;
                signal d1_jtag_uart_avalon_jtag_slave_end_xfer :  STD_LOGIC;
                signal d1_lcd_display_control_slave_end_xfer :  STD_LOGIC;
                signal d1_led_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_packet_memory_s1_end_xfer :  STD_LOGIC;
                signal d1_packet_memory_s2_end_xfer :  STD_LOGIC;
                signal d1_pipeline_bridge_s1_end_xfer :  STD_LOGIC;
                signal d1_pll_s1_end_xfer :  STD_LOGIC;
                signal d1_reconfig_request_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_seven_seg_pio_s1_end_xfer :  STD_LOGIC;
                signal d1_sgdma_rx_csr_end_xfer :  STD_LOGIC;
                signal d1_sgdma_tx_csr_end_xfer :  STD_LOGIC;
                signal d1_sys_clk_timer_s1_end_xfer :  STD_LOGIC;
                signal d1_tse_mac_control_port_end_xfer :  STD_LOGIC;
                signal d1_tse_pll_s1_end_xfer :  STD_LOGIC;
                signal d1_uart1_s1_end_xfer :  STD_LOGIC;
                signal ddr_sdram_0_s1_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal ddr_sdram_0_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal ddr_sdram_0_s1_read :  STD_LOGIC;
                signal ddr_sdram_0_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ddr_sdram_0_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ddr_sdram_0_s1_readdatavalid :  STD_LOGIC;
                signal ddr_sdram_0_s1_reset_n :  STD_LOGIC;
                signal ddr_sdram_0_s1_waitrequest_n :  STD_LOGIC;
                signal ddr_sdram_0_s1_waitrequest_n_from_sa :  STD_LOGIC;
                signal ddr_sdram_0_s1_write :  STD_LOGIC;
                signal ddr_sdram_0_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal descriptor_memory_s1_address :  STD_LOGIC_VECTOR (10 DOWNTO 0);
                signal descriptor_memory_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal descriptor_memory_s1_chipselect :  STD_LOGIC;
                signal descriptor_memory_s1_clken :  STD_LOGIC;
                signal descriptor_memory_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal descriptor_memory_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal descriptor_memory_s1_write :  STD_LOGIC;
                signal descriptor_memory_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal ext_flash_s1_wait_counter_eq_0 :  STD_LOGIC;
                signal high_res_timer_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal high_res_timer_s1_chipselect :  STD_LOGIC;
                signal high_res_timer_s1_irq :  STD_LOGIC;
                signal high_res_timer_s1_irq_from_sa :  STD_LOGIC;
                signal high_res_timer_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal high_res_timer_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal high_res_timer_s1_reset_n :  STD_LOGIC;
                signal high_res_timer_s1_write_n :  STD_LOGIC;
                signal high_res_timer_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal incoming_ext_ssram_bus_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal internal_LCD_E_from_the_lcd_display :  STD_LOGIC;
                signal internal_LCD_RS_from_the_lcd_display :  STD_LOGIC;
                signal internal_LCD_RW_from_the_lcd_display :  STD_LOGIC;
                signal internal_adsc_n_to_the_ext_ssram :  STD_LOGIC;
                signal internal_bw_n_to_the_ext_ssram :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_bwe_n_to_the_ext_ssram :  STD_LOGIC;
                signal internal_chipenable1_n_to_the_ext_ssram :  STD_LOGIC;
                signal internal_clk_to_sdram_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal internal_clk_to_sdram_n_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal internal_ddr_a_from_the_ddr_sdram_0 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal internal_ddr_ba_from_the_ddr_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_ddr_cas_n_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal internal_ddr_cke_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal internal_ddr_cs_n_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal internal_ddr_dm_from_the_ddr_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal internal_ddr_ras_n_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal internal_ddr_we_n_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal internal_ena_10_from_the_tse_mac :  STD_LOGIC;
                signal internal_eth_mode_from_the_tse_mac :  STD_LOGIC;
                signal internal_ext_flash_enet_bus_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal internal_ext_ssram_bus_address :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal internal_gm_tx_d_from_the_tse_mac :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_gm_tx_en_from_the_tse_mac :  STD_LOGIC;
                signal internal_gm_tx_err_from_the_tse_mac :  STD_LOGIC;
                signal internal_jtag_debug_offchip_trace_clk_from_the_cpu :  STD_LOGIC;
                signal internal_jtag_debug_offchip_trace_data_from_the_cpu :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal internal_jtag_debug_trigout_from_the_cpu :  STD_LOGIC;
                signal internal_m_tx_d_from_the_tse_mac :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal internal_m_tx_en_from_the_tse_mac :  STD_LOGIC;
                signal internal_m_tx_err_from_the_tse_mac :  STD_LOGIC;
                signal internal_mdc_from_the_tse_mac :  STD_LOGIC;
                signal internal_mdio_oen_from_the_tse_mac :  STD_LOGIC;
                signal internal_mdio_out_from_the_tse_mac :  STD_LOGIC;
                signal internal_out_port_from_the_led_pio :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal internal_out_port_from_the_seven_seg_pio :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal internal_outputenable_n_to_the_ext_ssram :  STD_LOGIC;
                signal internal_pll_c0_out :  STD_LOGIC;
                signal internal_read_n_to_the_ext_flash :  STD_LOGIC;
                signal internal_select_n_to_the_ext_flash :  STD_LOGIC;
                signal internal_stratix_dll_control_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal internal_txd_from_the_uart1 :  STD_LOGIC;
                signal internal_write_n_to_the_ext_flash :  STD_LOGIC;
                signal interrupt_vector_interrupt_vector_estatus :  STD_LOGIC;
                signal interrupt_vector_interrupt_vector_ipending :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal interrupt_vector_interrupt_vector_result :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal interrupt_vector_interrupt_vector_result_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal interrupt_vector_interrupt_vector_select :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_address :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_chipselect :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_irq_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_read_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal jtag_uart_avalon_jtag_slave_readyfordata :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_reset_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_waitrequest_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_write_n :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal lcd_display_control_slave_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal lcd_display_control_slave_begintransfer :  STD_LOGIC;
                signal lcd_display_control_slave_read :  STD_LOGIC;
                signal lcd_display_control_slave_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal lcd_display_control_slave_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal lcd_display_control_slave_wait_counter_eq_0 :  STD_LOGIC;
                signal lcd_display_control_slave_write :  STD_LOGIC;
                signal lcd_display_control_slave_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal led_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal led_pio_s1_chipselect :  STD_LOGIC;
                signal led_pio_s1_readdata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal led_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal led_pio_s1_reset_n :  STD_LOGIC;
                signal led_pio_s1_write_n :  STD_LOGIC;
                signal led_pio_s1_writedata :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal module_input15 :  STD_LOGIC;
                signal module_input16 :  STD_LOGIC;
                signal module_input17 :  STD_LOGIC;
                signal out_clk_pll_c0 :  STD_LOGIC;
                signal out_clk_pll_c1 :  STD_LOGIC;
                signal out_clk_pll_c2 :  STD_LOGIC;
                signal out_clk_tse_pll_c0 :  STD_LOGIC;
                signal packet_memory_s1_address :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal packet_memory_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal packet_memory_s1_chipselect :  STD_LOGIC;
                signal packet_memory_s1_clken :  STD_LOGIC;
                signal packet_memory_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal packet_memory_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal packet_memory_s1_write :  STD_LOGIC;
                signal packet_memory_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal packet_memory_s2_address :  STD_LOGIC_VECTOR (13 DOWNTO 0);
                signal packet_memory_s2_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal packet_memory_s2_chipselect :  STD_LOGIC;
                signal packet_memory_s2_clken :  STD_LOGIC;
                signal packet_memory_s2_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal packet_memory_s2_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal packet_memory_s2_write :  STD_LOGIC;
                signal packet_memory_s2_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pipeline_bridge_m1_address :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pipeline_bridge_m1_address_to_slave :  STD_LOGIC_VECTOR (24 DOWNTO 0);
                signal pipeline_bridge_m1_burstcount :  STD_LOGIC;
                signal pipeline_bridge_m1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pipeline_bridge_m1_byteenable_ext_flash_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_chipselect :  STD_LOGIC;
                signal pipeline_bridge_m1_dbs_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_m1_dbs_write_8 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal pipeline_bridge_m1_debugaccess :  STD_LOGIC;
                signal pipeline_bridge_m1_endofpacket :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_button_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_cpu_jtag_debug_module :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_ext_flash_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_high_res_timer_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_lcd_display_control_slave :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_led_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_reconfig_request_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_seven_seg_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_sgdma_rx_csr :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_sgdma_tx_csr :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_sys_clk_timer_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_granted_uart1_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_latency_counter :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_button_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_ext_flash_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_high_res_timer_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_lcd_display_control_slave :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_led_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_sgdma_rx_csr :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_sgdma_tx_csr :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_qualified_request_uart1_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_read :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_button_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_ext_flash_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_high_res_timer_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_lcd_display_control_slave :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_led_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_sgdma_rx_csr :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_sgdma_tx_csr :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_read_data_valid_uart1_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pipeline_bridge_m1_readdatavalid :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_button_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_cpu_jtag_debug_module :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_ext_flash_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_high_res_timer_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_lcd_display_control_slave :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_led_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_reconfig_request_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_seven_seg_pio_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_sgdma_rx_csr :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_sgdma_tx_csr :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_sys_clk_timer_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_requests_uart1_s1 :  STD_LOGIC;
                signal pipeline_bridge_m1_waitrequest :  STD_LOGIC;
                signal pipeline_bridge_m1_write :  STD_LOGIC;
                signal pipeline_bridge_m1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pipeline_bridge_s1_address :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal pipeline_bridge_s1_arbiterlock :  STD_LOGIC;
                signal pipeline_bridge_s1_arbiterlock2 :  STD_LOGIC;
                signal pipeline_bridge_s1_burstcount :  STD_LOGIC;
                signal pipeline_bridge_s1_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal pipeline_bridge_s1_chipselect :  STD_LOGIC;
                signal pipeline_bridge_s1_debugaccess :  STD_LOGIC;
                signal pipeline_bridge_s1_endofpacket :  STD_LOGIC;
                signal pipeline_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal pipeline_bridge_s1_nativeaddress :  STD_LOGIC_VECTOR (22 DOWNTO 0);
                signal pipeline_bridge_s1_read :  STD_LOGIC;
                signal pipeline_bridge_s1_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pipeline_bridge_s1_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pipeline_bridge_s1_readdatavalid :  STD_LOGIC;
                signal pipeline_bridge_s1_reset_n :  STD_LOGIC;
                signal pipeline_bridge_s1_waitrequest :  STD_LOGIC;
                signal pipeline_bridge_s1_waitrequest_from_sa :  STD_LOGIC;
                signal pipeline_bridge_s1_write :  STD_LOGIC;
                signal pipeline_bridge_s1_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal pll_c0_out_reset_n :  STD_LOGIC;
                signal pll_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal pll_s1_chipselect :  STD_LOGIC;
                signal pll_s1_read :  STD_LOGIC;
                signal pll_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pll_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal pll_s1_reset_n :  STD_LOGIC;
                signal pll_s1_resetrequest :  STD_LOGIC;
                signal pll_s1_resetrequest_from_sa :  STD_LOGIC;
                signal pll_s1_write :  STD_LOGIC;
                signal pll_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal reconfig_request_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal reconfig_request_pio_s1_chipselect :  STD_LOGIC;
                signal reconfig_request_pio_s1_readdata :  STD_LOGIC;
                signal reconfig_request_pio_s1_readdata_from_sa :  STD_LOGIC;
                signal reconfig_request_pio_s1_reset_n :  STD_LOGIC;
                signal reconfig_request_pio_s1_write_n :  STD_LOGIC;
                signal reconfig_request_pio_s1_writedata :  STD_LOGIC;
                signal reset_n_sources :  STD_LOGIC;
                signal seven_seg_pio_s1_address :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal seven_seg_pio_s1_chipselect :  STD_LOGIC;
                signal seven_seg_pio_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal seven_seg_pio_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal seven_seg_pio_s1_reset_n :  STD_LOGIC;
                signal seven_seg_pio_s1_write_n :  STD_LOGIC;
                signal seven_seg_pio_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sgdma_rx_csr_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal sgdma_rx_csr_chipselect :  STD_LOGIC;
                signal sgdma_rx_csr_irq :  STD_LOGIC;
                signal sgdma_rx_csr_irq_from_sa :  STD_LOGIC;
                signal sgdma_rx_csr_read :  STD_LOGIC;
                signal sgdma_rx_csr_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_csr_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_csr_reset_n :  STD_LOGIC;
                signal sgdma_rx_csr_write :  STD_LOGIC;
                signal sgdma_rx_csr_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_read_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_read_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_latency_counter :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_read_readdatavalid :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_read_waitrequest :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_descriptor_write_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_waitrequest :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_write :  STD_LOGIC;
                signal sgdma_rx_descriptor_write_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_in_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_in_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sgdma_rx_in_endofpacket :  STD_LOGIC;
                signal sgdma_rx_in_error :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal sgdma_rx_in_ready :  STD_LOGIC;
                signal sgdma_rx_in_ready_from_sa :  STD_LOGIC;
                signal sgdma_rx_in_startofpacket :  STD_LOGIC;
                signal sgdma_rx_in_valid :  STD_LOGIC;
                signal sgdma_rx_m_write_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_m_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_rx_m_write_byteenable :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal sgdma_rx_m_write_granted_ddr_sdram_0_s1 :  STD_LOGIC;
                signal sgdma_rx_m_write_granted_ext_ssram_s1 :  STD_LOGIC;
                signal sgdma_rx_m_write_granted_packet_memory_s2 :  STD_LOGIC;
                signal sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 :  STD_LOGIC;
                signal sgdma_rx_m_write_qualified_request_ext_ssram_s1 :  STD_LOGIC;
                signal sgdma_rx_m_write_qualified_request_packet_memory_s2 :  STD_LOGIC;
                signal sgdma_rx_m_write_requests_ddr_sdram_0_s1 :  STD_LOGIC;
                signal sgdma_rx_m_write_requests_ext_ssram_s1 :  STD_LOGIC;
                signal sgdma_rx_m_write_requests_packet_memory_s2 :  STD_LOGIC;
                signal sgdma_rx_m_write_waitrequest :  STD_LOGIC;
                signal sgdma_rx_m_write_write :  STD_LOGIC;
                signal sgdma_rx_m_write_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_csr_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal sgdma_tx_csr_chipselect :  STD_LOGIC;
                signal sgdma_tx_csr_irq :  STD_LOGIC;
                signal sgdma_tx_csr_irq_from_sa :  STD_LOGIC;
                signal sgdma_tx_csr_read :  STD_LOGIC;
                signal sgdma_tx_csr_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_csr_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_csr_reset_n :  STD_LOGIC;
                signal sgdma_tx_csr_write :  STD_LOGIC;
                signal sgdma_tx_csr_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_read_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_read_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_latency_counter :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_read_readdatavalid :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_read_waitrequest :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_write_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_descriptor_write_granted_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_requests_descriptor_memory_s1 :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_waitrequest :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_write :  STD_LOGIC;
                signal sgdma_tx_descriptor_write_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_m_read_address :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_m_read_address_to_slave :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_m_read_granted_ddr_sdram_0_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_granted_ext_ssram_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_granted_packet_memory_s2 :  STD_LOGIC;
                signal sgdma_tx_m_read_latency_counter :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_qualified_request_ext_ssram_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_qualified_request_packet_memory_s2 :  STD_LOGIC;
                signal sgdma_tx_m_read_read :  STD_LOGIC;
                signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register :  STD_LOGIC;
                signal sgdma_tx_m_read_read_data_valid_ext_ssram_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_read_data_valid_packet_memory_s2 :  STD_LOGIC;
                signal sgdma_tx_m_read_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_m_read_readdatavalid :  STD_LOGIC;
                signal sgdma_tx_m_read_requests_ddr_sdram_0_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_requests_ext_ssram_s1 :  STD_LOGIC;
                signal sgdma_tx_m_read_requests_packet_memory_s2 :  STD_LOGIC;
                signal sgdma_tx_m_read_waitrequest :  STD_LOGIC;
                signal sgdma_tx_out_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal sgdma_tx_out_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal sgdma_tx_out_endofpacket :  STD_LOGIC;
                signal sgdma_tx_out_error :  STD_LOGIC;
                signal sgdma_tx_out_ready :  STD_LOGIC;
                signal sgdma_tx_out_startofpacket :  STD_LOGIC;
                signal sgdma_tx_out_valid :  STD_LOGIC;
                signal sys_clk_timer_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal sys_clk_timer_s1_chipselect :  STD_LOGIC;
                signal sys_clk_timer_s1_irq :  STD_LOGIC;
                signal sys_clk_timer_s1_irq_from_sa :  STD_LOGIC;
                signal sys_clk_timer_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sys_clk_timer_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal sys_clk_timer_s1_reset_n :  STD_LOGIC;
                signal sys_clk_timer_s1_write_n :  STD_LOGIC;
                signal sys_clk_timer_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal tse_mac_control_port_address :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal tse_mac_control_port_read :  STD_LOGIC;
                signal tse_mac_control_port_readdata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_control_port_readdata_from_sa :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_control_port_reset :  STD_LOGIC;
                signal tse_mac_control_port_waitrequest :  STD_LOGIC;
                signal tse_mac_control_port_waitrequest_from_sa :  STD_LOGIC;
                signal tse_mac_control_port_write :  STD_LOGIC;
                signal tse_mac_control_port_writedata :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_receive_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_receive_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tse_mac_receive_endofpacket :  STD_LOGIC;
                signal tse_mac_receive_error :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal tse_mac_receive_ready :  STD_LOGIC;
                signal tse_mac_receive_startofpacket :  STD_LOGIC;
                signal tse_mac_receive_valid :  STD_LOGIC;
                signal tse_mac_transmit_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal tse_mac_transmit_empty :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal tse_mac_transmit_endofpacket :  STD_LOGIC;
                signal tse_mac_transmit_error :  STD_LOGIC;
                signal tse_mac_transmit_ready :  STD_LOGIC;
                signal tse_mac_transmit_ready_from_sa :  STD_LOGIC;
                signal tse_mac_transmit_startofpacket :  STD_LOGIC;
                signal tse_mac_transmit_valid :  STD_LOGIC;
                signal tse_pll_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal tse_pll_s1_chipselect :  STD_LOGIC;
                signal tse_pll_s1_read :  STD_LOGIC;
                signal tse_pll_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal tse_pll_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal tse_pll_s1_reset_n :  STD_LOGIC;
                signal tse_pll_s1_resetrequest :  STD_LOGIC;
                signal tse_pll_s1_resetrequest_from_sa :  STD_LOGIC;
                signal tse_pll_s1_write :  STD_LOGIC;
                signal tse_pll_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal uart1_s1_address :  STD_LOGIC_VECTOR (2 DOWNTO 0);
                signal uart1_s1_begintransfer :  STD_LOGIC;
                signal uart1_s1_chipselect :  STD_LOGIC;
                signal uart1_s1_dataavailable :  STD_LOGIC;
                signal uart1_s1_dataavailable_from_sa :  STD_LOGIC;
                signal uart1_s1_irq :  STD_LOGIC;
                signal uart1_s1_irq_from_sa :  STD_LOGIC;
                signal uart1_s1_read_n :  STD_LOGIC;
                signal uart1_s1_readdata :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal uart1_s1_readdata_from_sa :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal uart1_s1_readyfordata :  STD_LOGIC;
                signal uart1_s1_readyfordata_from_sa :  STD_LOGIC;
                signal uart1_s1_reset_n :  STD_LOGIC;
                signal uart1_s1_write_n :  STD_LOGIC;
                signal uart1_s1_writedata :  STD_LOGIC_VECTOR (15 DOWNTO 0);

begin

  --the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in, which is an e_instance
  the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_arbitrator
    port map(
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_address => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_address,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_byteenable => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_byteenable,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_nativeaddress => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_nativeaddress,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_read => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_read,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reset_n => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reset_n,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_write => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_write,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_writedata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_writedata,
      d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer => d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer,
      pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in => pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in,
      pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in => pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in,
      pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in => pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in,
      pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in => pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest,
      clk => internal_pll_c0_out,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_byteenable => pipeline_bridge_m1_byteenable,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n
    );


  --the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out, which is an e_instance
  the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_arbitrator
    port map(
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_readdata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_readdata,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_reset_n => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_reset_n,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_data_valid_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_data_valid_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata,
      clk => clk,
      d1_pll_s1_end_xfer => d1_pll_s1_end_xfer,
      pll_s1_readdata_from_sa => pll_s1_readdata_from_sa,
      reset_n => clk_reset_n
    );


  --the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0, which is an e_ptf_instance
  the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0 : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0
    port map(
      master_address => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address,
      master_byteenable => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_byteenable,
      master_nativeaddress => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_nativeaddress,
      master_read => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read,
      master_write => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write,
      master_writedata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata,
      slave_endofpacket => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket,
      slave_readdata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata,
      slave_waitrequest => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest,
      master_clk => clk,
      master_endofpacket => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_endofpacket,
      master_readdata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_readdata,
      master_reset_n => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_reset_n,
      master_waitrequest => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_waitrequest,
      slave_address => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_address,
      slave_byteenable => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_byteenable,
      slave_clk => internal_pll_c0_out,
      slave_nativeaddress => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_nativeaddress,
      slave_read => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_read,
      slave_reset_n => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_reset_n,
      slave_write => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_write,
      slave_writedata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_writedata
    );


  --the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in, which is an e_instance
  the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_arbitrator
    port map(
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_address => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_address,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_byteenable => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_byteenable,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_nativeaddress => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_nativeaddress,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_read => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_read,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reset_n => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reset_n,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_write => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_write,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_writedata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_writedata,
      d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer => d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer,
      pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in => pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in,
      pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in => pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in,
      pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in => pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in,
      pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in => pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest,
      clk => internal_pll_c0_out,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_byteenable => pipeline_bridge_m1_byteenable,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n
    );


  --the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out, which is an e_instance
  the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_arbitrator
    port map(
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_readdata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_readdata,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_reset_n => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_reset_n,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_data_valid_tse_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_data_valid_tse_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata,
      clk => clk_to_tse_pll,
      d1_tse_pll_s1_end_xfer => d1_tse_pll_s1_end_xfer,
      reset_n => clk_to_tse_pll_reset_n,
      tse_pll_s1_readdata_from_sa => tse_pll_s1_readdata_from_sa
    );


  --the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1, which is an e_ptf_instance
  the_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1 : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1
    port map(
      master_address => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address,
      master_byteenable => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_byteenable,
      master_nativeaddress => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_nativeaddress,
      master_read => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read,
      master_write => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write,
      master_writedata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata,
      slave_endofpacket => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket,
      slave_readdata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata,
      slave_waitrequest => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest,
      master_clk => clk_to_tse_pll,
      master_endofpacket => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_endofpacket,
      master_readdata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_readdata,
      master_reset_n => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_reset_n,
      master_waitrequest => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_waitrequest,
      slave_address => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_address,
      slave_byteenable => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_byteenable,
      slave_clk => internal_pll_c0_out,
      slave_nativeaddress => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_nativeaddress,
      slave_read => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_read,
      slave_reset_n => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_reset_n,
      slave_write => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_write,
      slave_writedata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_writedata
    );


  --the_bswap_s1, which is an e_instance
  the_bswap_s1 : bswap_s1_arbitrator
    port map(
      bswap_s1_dataa => bswap_s1_dataa,
      bswap_s1_datab => bswap_s1_datab,
      bswap_s1_result_from_sa => bswap_s1_result_from_sa,
      bswap_s1_result => bswap_s1_result,
      bswap_s1_select => bswap_s1_select,
      clk => internal_pll_c0_out,
      cpu_custom_instruction_master_combo_dataa => cpu_custom_instruction_master_combo_dataa,
      cpu_custom_instruction_master_combo_datab => cpu_custom_instruction_master_combo_datab,
      reset_n => pll_c0_out_reset_n
    );


  --the_bswap, which is an e_ptf_instance
  the_bswap : bswap
    port map(
      result => bswap_s1_result,
      dataa => bswap_s1_dataa,
      datab => bswap_s1_datab
    );


  --the_button_pio_s1, which is an e_instance
  the_button_pio_s1 : button_pio_s1_arbitrator
    port map(
      button_pio_s1_address => button_pio_s1_address,
      button_pio_s1_chipselect => button_pio_s1_chipselect,
      button_pio_s1_irq_from_sa => button_pio_s1_irq_from_sa,
      button_pio_s1_readdata_from_sa => button_pio_s1_readdata_from_sa,
      button_pio_s1_reset_n => button_pio_s1_reset_n,
      button_pio_s1_write_n => button_pio_s1_write_n,
      button_pio_s1_writedata => button_pio_s1_writedata,
      d1_button_pio_s1_end_xfer => d1_button_pio_s1_end_xfer,
      pipeline_bridge_m1_granted_button_pio_s1 => pipeline_bridge_m1_granted_button_pio_s1,
      pipeline_bridge_m1_qualified_request_button_pio_s1 => pipeline_bridge_m1_qualified_request_button_pio_s1,
      pipeline_bridge_m1_read_data_valid_button_pio_s1 => pipeline_bridge_m1_read_data_valid_button_pio_s1,
      pipeline_bridge_m1_requests_button_pio_s1 => pipeline_bridge_m1_requests_button_pio_s1,
      button_pio_s1_irq => button_pio_s1_irq,
      button_pio_s1_readdata => button_pio_s1_readdata,
      clk => internal_pll_c0_out,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n
    );


  --the_button_pio, which is an e_ptf_instance
  the_button_pio : button_pio
    port map(
      irq => button_pio_s1_irq,
      readdata => button_pio_s1_readdata,
      address => button_pio_s1_address,
      chipselect => button_pio_s1_chipselect,
      clk => internal_pll_c0_out,
      in_port => in_port_to_the_button_pio,
      reset_n => button_pio_s1_reset_n,
      write_n => button_pio_s1_write_n,
      writedata => button_pio_s1_writedata
    );


  --the_cpu_jtag_debug_module, which is an e_instance
  the_cpu_jtag_debug_module : cpu_jtag_debug_module_arbitrator
    port map(
      cpu_jtag_debug_module_address => cpu_jtag_debug_module_address,
      cpu_jtag_debug_module_begintransfer => cpu_jtag_debug_module_begintransfer,
      cpu_jtag_debug_module_byteenable => cpu_jtag_debug_module_byteenable,
      cpu_jtag_debug_module_chipselect => cpu_jtag_debug_module_chipselect,
      cpu_jtag_debug_module_debugaccess => cpu_jtag_debug_module_debugaccess,
      cpu_jtag_debug_module_readdata_from_sa => cpu_jtag_debug_module_readdata_from_sa,
      cpu_jtag_debug_module_reset => cpu_jtag_debug_module_reset,
      cpu_jtag_debug_module_resetrequest_from_sa => cpu_jtag_debug_module_resetrequest_from_sa,
      cpu_jtag_debug_module_write => cpu_jtag_debug_module_write,
      cpu_jtag_debug_module_writedata => cpu_jtag_debug_module_writedata,
      d1_cpu_jtag_debug_module_end_xfer => d1_cpu_jtag_debug_module_end_xfer,
      pipeline_bridge_m1_granted_cpu_jtag_debug_module => pipeline_bridge_m1_granted_cpu_jtag_debug_module,
      pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module => pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module,
      pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module => pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module,
      pipeline_bridge_m1_requests_cpu_jtag_debug_module => pipeline_bridge_m1_requests_cpu_jtag_debug_module,
      clk => internal_pll_c0_out,
      cpu_jtag_debug_module_readdata => cpu_jtag_debug_module_readdata,
      cpu_jtag_debug_module_resetrequest => cpu_jtag_debug_module_resetrequest,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_byteenable => pipeline_bridge_m1_byteenable,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_debugaccess => pipeline_bridge_m1_debugaccess,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n
    );


  --the_cpu_custom_instruction_master, which is an e_instance
  the_cpu_custom_instruction_master : cpu_custom_instruction_master_arbitrator
    port map(
      bswap_s1_select => bswap_s1_select,
      cpu_custom_instruction_master_combo_result => cpu_custom_instruction_master_combo_result,
      cpu_custom_instruction_master_reset_n => cpu_custom_instruction_master_reset_n,
      interrupt_vector_interrupt_vector_select => interrupt_vector_interrupt_vector_select,
      bswap_s1_result_from_sa => bswap_s1_result_from_sa,
      clk => internal_pll_c0_out,
      cpu_custom_instruction_master_combo_n => cpu_custom_instruction_master_combo_n,
      interrupt_vector_interrupt_vector_result_from_sa => interrupt_vector_interrupt_vector_result_from_sa,
      reset_n => pll_c0_out_reset_n
    );


  --the_cpu_data_master, which is an e_instance
  the_cpu_data_master : cpu_data_master_arbitrator
    port map(
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_irq => cpu_data_master_irq,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_readdata => cpu_data_master_readdata,
      cpu_data_master_readdatavalid => cpu_data_master_readdatavalid,
      cpu_data_master_waitrequest => cpu_data_master_waitrequest,
      button_pio_s1_irq_from_sa => button_pio_s1_irq_from_sa,
      clk => internal_pll_c0_out,
      cpu_data_master_address => cpu_data_master_address,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_granted_ddr_sdram_0_s1 => cpu_data_master_granted_ddr_sdram_0_s1,
      cpu_data_master_granted_descriptor_memory_s1 => cpu_data_master_granted_descriptor_memory_s1,
      cpu_data_master_granted_ext_ssram_s1 => cpu_data_master_granted_ext_ssram_s1,
      cpu_data_master_granted_packet_memory_s1 => cpu_data_master_granted_packet_memory_s1,
      cpu_data_master_granted_pipeline_bridge_s1 => cpu_data_master_granted_pipeline_bridge_s1,
      cpu_data_master_granted_tse_mac_control_port => cpu_data_master_granted_tse_mac_control_port,
      cpu_data_master_qualified_request_ddr_sdram_0_s1 => cpu_data_master_qualified_request_ddr_sdram_0_s1,
      cpu_data_master_qualified_request_descriptor_memory_s1 => cpu_data_master_qualified_request_descriptor_memory_s1,
      cpu_data_master_qualified_request_ext_ssram_s1 => cpu_data_master_qualified_request_ext_ssram_s1,
      cpu_data_master_qualified_request_packet_memory_s1 => cpu_data_master_qualified_request_packet_memory_s1,
      cpu_data_master_qualified_request_pipeline_bridge_s1 => cpu_data_master_qualified_request_pipeline_bridge_s1,
      cpu_data_master_qualified_request_tse_mac_control_port => cpu_data_master_qualified_request_tse_mac_control_port,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_ddr_sdram_0_s1 => cpu_data_master_read_data_valid_ddr_sdram_0_s1,
      cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      cpu_data_master_read_data_valid_descriptor_memory_s1 => cpu_data_master_read_data_valid_descriptor_memory_s1,
      cpu_data_master_read_data_valid_ext_ssram_s1 => cpu_data_master_read_data_valid_ext_ssram_s1,
      cpu_data_master_read_data_valid_packet_memory_s1 => cpu_data_master_read_data_valid_packet_memory_s1,
      cpu_data_master_read_data_valid_pipeline_bridge_s1 => cpu_data_master_read_data_valid_pipeline_bridge_s1,
      cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register,
      cpu_data_master_read_data_valid_tse_mac_control_port => cpu_data_master_read_data_valid_tse_mac_control_port,
      cpu_data_master_requests_ddr_sdram_0_s1 => cpu_data_master_requests_ddr_sdram_0_s1,
      cpu_data_master_requests_descriptor_memory_s1 => cpu_data_master_requests_descriptor_memory_s1,
      cpu_data_master_requests_ext_ssram_s1 => cpu_data_master_requests_ext_ssram_s1,
      cpu_data_master_requests_packet_memory_s1 => cpu_data_master_requests_packet_memory_s1,
      cpu_data_master_requests_pipeline_bridge_s1 => cpu_data_master_requests_pipeline_bridge_s1,
      cpu_data_master_requests_tse_mac_control_port => cpu_data_master_requests_tse_mac_control_port,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      d1_ddr_sdram_0_s1_end_xfer => d1_ddr_sdram_0_s1_end_xfer,
      d1_descriptor_memory_s1_end_xfer => d1_descriptor_memory_s1_end_xfer,
      d1_ext_ssram_bus_avalon_slave_end_xfer => d1_ext_ssram_bus_avalon_slave_end_xfer,
      d1_packet_memory_s1_end_xfer => d1_packet_memory_s1_end_xfer,
      d1_pipeline_bridge_s1_end_xfer => d1_pipeline_bridge_s1_end_xfer,
      d1_tse_mac_control_port_end_xfer => d1_tse_mac_control_port_end_xfer,
      ddr_sdram_0_s1_readdata_from_sa => ddr_sdram_0_s1_readdata_from_sa,
      ddr_sdram_0_s1_waitrequest_n_from_sa => ddr_sdram_0_s1_waitrequest_n_from_sa,
      descriptor_memory_s1_readdata_from_sa => descriptor_memory_s1_readdata_from_sa,
      high_res_timer_s1_irq_from_sa => high_res_timer_s1_irq_from_sa,
      incoming_ext_ssram_bus_data => incoming_ext_ssram_bus_data,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      packet_memory_s1_readdata_from_sa => packet_memory_s1_readdata_from_sa,
      pipeline_bridge_s1_readdata_from_sa => pipeline_bridge_s1_readdata_from_sa,
      pipeline_bridge_s1_waitrequest_from_sa => pipeline_bridge_s1_waitrequest_from_sa,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_csr_irq_from_sa => sgdma_rx_csr_irq_from_sa,
      sgdma_tx_csr_irq_from_sa => sgdma_tx_csr_irq_from_sa,
      sys_clk_timer_s1_irq_from_sa => sys_clk_timer_s1_irq_from_sa,
      tse_mac_control_port_readdata_from_sa => tse_mac_control_port_readdata_from_sa,
      tse_mac_control_port_waitrequest_from_sa => tse_mac_control_port_waitrequest_from_sa,
      uart1_s1_irq_from_sa => uart1_s1_irq_from_sa
    );


  --the_cpu_instruction_master, which is an e_instance
  the_cpu_instruction_master : cpu_instruction_master_arbitrator
    port map(
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_readdata => cpu_instruction_master_readdata,
      cpu_instruction_master_readdatavalid => cpu_instruction_master_readdatavalid,
      cpu_instruction_master_waitrequest => cpu_instruction_master_waitrequest,
      clk => internal_pll_c0_out,
      cpu_instruction_master_address => cpu_instruction_master_address,
      cpu_instruction_master_granted_ddr_sdram_0_s1 => cpu_instruction_master_granted_ddr_sdram_0_s1,
      cpu_instruction_master_granted_ext_ssram_s1 => cpu_instruction_master_granted_ext_ssram_s1,
      cpu_instruction_master_granted_pipeline_bridge_s1 => cpu_instruction_master_granted_pipeline_bridge_s1,
      cpu_instruction_master_qualified_request_ddr_sdram_0_s1 => cpu_instruction_master_qualified_request_ddr_sdram_0_s1,
      cpu_instruction_master_qualified_request_ext_ssram_s1 => cpu_instruction_master_qualified_request_ext_ssram_s1,
      cpu_instruction_master_qualified_request_pipeline_bridge_s1 => cpu_instruction_master_qualified_request_pipeline_bridge_s1,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_ddr_sdram_0_s1 => cpu_instruction_master_read_data_valid_ddr_sdram_0_s1,
      cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      cpu_instruction_master_read_data_valid_ext_ssram_s1 => cpu_instruction_master_read_data_valid_ext_ssram_s1,
      cpu_instruction_master_read_data_valid_pipeline_bridge_s1 => cpu_instruction_master_read_data_valid_pipeline_bridge_s1,
      cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register,
      cpu_instruction_master_requests_ddr_sdram_0_s1 => cpu_instruction_master_requests_ddr_sdram_0_s1,
      cpu_instruction_master_requests_ext_ssram_s1 => cpu_instruction_master_requests_ext_ssram_s1,
      cpu_instruction_master_requests_pipeline_bridge_s1 => cpu_instruction_master_requests_pipeline_bridge_s1,
      d1_ddr_sdram_0_s1_end_xfer => d1_ddr_sdram_0_s1_end_xfer,
      d1_ext_ssram_bus_avalon_slave_end_xfer => d1_ext_ssram_bus_avalon_slave_end_xfer,
      d1_pipeline_bridge_s1_end_xfer => d1_pipeline_bridge_s1_end_xfer,
      ddr_sdram_0_s1_readdata_from_sa => ddr_sdram_0_s1_readdata_from_sa,
      ddr_sdram_0_s1_waitrequest_n_from_sa => ddr_sdram_0_s1_waitrequest_n_from_sa,
      incoming_ext_ssram_bus_data => incoming_ext_ssram_bus_data,
      pipeline_bridge_s1_readdata_from_sa => pipeline_bridge_s1_readdata_from_sa,
      pipeline_bridge_s1_waitrequest_from_sa => pipeline_bridge_s1_waitrequest_from_sa,
      reset_n => pll_c0_out_reset_n
    );


  --the_cpu, which is an e_ptf_instance
  the_cpu : cpu
    port map(
      E_ci_combo_a => cpu_custom_instruction_master_combo_a,
      E_ci_combo_b => cpu_custom_instruction_master_combo_b,
      E_ci_combo_c => cpu_custom_instruction_master_combo_c,
      E_ci_combo_dataa => cpu_custom_instruction_master_combo_dataa,
      E_ci_combo_datab => cpu_custom_instruction_master_combo_datab,
      E_ci_combo_estatus => cpu_custom_instruction_master_combo_estatus,
      E_ci_combo_ipending => cpu_custom_instruction_master_combo_ipending,
      E_ci_combo_n => cpu_custom_instruction_master_combo_n,
      E_ci_combo_readra => cpu_custom_instruction_master_combo_readra,
      E_ci_combo_readrb => cpu_custom_instruction_master_combo_readrb,
      E_ci_combo_status => cpu_custom_instruction_master_combo_status,
      E_ci_combo_writerc => cpu_custom_instruction_master_combo_writerc,
      d_address => cpu_data_master_address,
      d_byteenable => cpu_data_master_byteenable,
      d_read => cpu_data_master_read,
      d_write => cpu_data_master_write,
      d_writedata => cpu_data_master_writedata,
      i_address => cpu_instruction_master_address,
      i_read => cpu_instruction_master_read,
      jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,
      jtag_debug_module_readdata => cpu_jtag_debug_module_readdata,
      jtag_debug_module_resetrequest => cpu_jtag_debug_module_resetrequest,
      jtag_debug_offchip_trace_clk => internal_jtag_debug_offchip_trace_clk_from_the_cpu,
      jtag_debug_offchip_trace_data => internal_jtag_debug_offchip_trace_data_from_the_cpu,
      jtag_debug_trigout => internal_jtag_debug_trigout_from_the_cpu,
      E_ci_combo_result => cpu_custom_instruction_master_combo_result,
      clk => internal_pll_c0_out,
      d_irq => cpu_data_master_irq,
      d_readdata => cpu_data_master_readdata,
      d_readdatavalid => cpu_data_master_readdatavalid,
      d_waitrequest => cpu_data_master_waitrequest,
      i_readdata => cpu_instruction_master_readdata,
      i_readdatavalid => cpu_instruction_master_readdatavalid,
      i_waitrequest => cpu_instruction_master_waitrequest,
      jtag_debug_module_address => cpu_jtag_debug_module_address,
      jtag_debug_module_begintransfer => cpu_jtag_debug_module_begintransfer,
      jtag_debug_module_byteenable => cpu_jtag_debug_module_byteenable,
      jtag_debug_module_clk => internal_pll_c0_out,
      jtag_debug_module_debugaccess => cpu_jtag_debug_module_debugaccess,
      jtag_debug_module_reset => cpu_jtag_debug_module_reset,
      jtag_debug_module_select => cpu_jtag_debug_module_chipselect,
      jtag_debug_module_write => cpu_jtag_debug_module_write,
      jtag_debug_module_writedata => cpu_jtag_debug_module_writedata,
      reset_n => cpu_custom_instruction_master_reset_n
    );


  --the_ddr_sdram_0_s1, which is an e_instance
  the_ddr_sdram_0_s1 : ddr_sdram_0_s1_arbitrator
    port map(
      cpu_data_master_granted_ddr_sdram_0_s1 => cpu_data_master_granted_ddr_sdram_0_s1,
      cpu_data_master_qualified_request_ddr_sdram_0_s1 => cpu_data_master_qualified_request_ddr_sdram_0_s1,
      cpu_data_master_read_data_valid_ddr_sdram_0_s1 => cpu_data_master_read_data_valid_ddr_sdram_0_s1,
      cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      cpu_data_master_requests_ddr_sdram_0_s1 => cpu_data_master_requests_ddr_sdram_0_s1,
      cpu_instruction_master_granted_ddr_sdram_0_s1 => cpu_instruction_master_granted_ddr_sdram_0_s1,
      cpu_instruction_master_qualified_request_ddr_sdram_0_s1 => cpu_instruction_master_qualified_request_ddr_sdram_0_s1,
      cpu_instruction_master_read_data_valid_ddr_sdram_0_s1 => cpu_instruction_master_read_data_valid_ddr_sdram_0_s1,
      cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      cpu_instruction_master_requests_ddr_sdram_0_s1 => cpu_instruction_master_requests_ddr_sdram_0_s1,
      d1_ddr_sdram_0_s1_end_xfer => d1_ddr_sdram_0_s1_end_xfer,
      ddr_sdram_0_s1_address => ddr_sdram_0_s1_address,
      ddr_sdram_0_s1_byteenable => ddr_sdram_0_s1_byteenable,
      ddr_sdram_0_s1_read => ddr_sdram_0_s1_read,
      ddr_sdram_0_s1_readdata_from_sa => ddr_sdram_0_s1_readdata_from_sa,
      ddr_sdram_0_s1_reset_n => ddr_sdram_0_s1_reset_n,
      ddr_sdram_0_s1_waitrequest_n_from_sa => ddr_sdram_0_s1_waitrequest_n_from_sa,
      ddr_sdram_0_s1_write => ddr_sdram_0_s1_write,
      ddr_sdram_0_s1_writedata => ddr_sdram_0_s1_writedata,
      sgdma_rx_m_write_granted_ddr_sdram_0_s1 => sgdma_rx_m_write_granted_ddr_sdram_0_s1,
      sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 => sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1,
      sgdma_rx_m_write_requests_ddr_sdram_0_s1 => sgdma_rx_m_write_requests_ddr_sdram_0_s1,
      sgdma_tx_m_read_granted_ddr_sdram_0_s1 => sgdma_tx_m_read_granted_ddr_sdram_0_s1,
      sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 => sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1,
      sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1 => sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1,
      sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register => sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register,
      sgdma_tx_m_read_requests_ddr_sdram_0_s1 => sgdma_tx_m_read_requests_ddr_sdram_0_s1,
      clk => internal_pll_c0_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register,
      ddr_sdram_0_s1_readdata => ddr_sdram_0_s1_readdata,
      ddr_sdram_0_s1_readdatavalid => ddr_sdram_0_s1_readdatavalid,
      ddr_sdram_0_s1_waitrequest_n => ddr_sdram_0_s1_waitrequest_n,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_m_write_address_to_slave => sgdma_rx_m_write_address_to_slave,
      sgdma_rx_m_write_byteenable => sgdma_rx_m_write_byteenable,
      sgdma_rx_m_write_write => sgdma_rx_m_write_write,
      sgdma_rx_m_write_writedata => sgdma_rx_m_write_writedata,
      sgdma_tx_m_read_address_to_slave => sgdma_tx_m_read_address_to_slave,
      sgdma_tx_m_read_latency_counter => sgdma_tx_m_read_latency_counter,
      sgdma_tx_m_read_read => sgdma_tx_m_read_read
    );


  --the_ddr_sdram_0, which is an e_ptf_instance
  the_ddr_sdram_0 : ddr_sdram_0
    port map(
      clk_to_sdram => internal_clk_to_sdram_from_the_ddr_sdram_0,
      clk_to_sdram_n => internal_clk_to_sdram_n_from_the_ddr_sdram_0,
      ddr_a => internal_ddr_a_from_the_ddr_sdram_0,
      ddr_ba => internal_ddr_ba_from_the_ddr_sdram_0,
      ddr_cas_n => internal_ddr_cas_n_from_the_ddr_sdram_0,
      ddr_cke => internal_ddr_cke_from_the_ddr_sdram_0,
      ddr_cs_n => internal_ddr_cs_n_from_the_ddr_sdram_0,
      ddr_dm => internal_ddr_dm_from_the_ddr_sdram_0,
      ddr_dq => ddr_dq_to_and_from_the_ddr_sdram_0,
      ddr_dqs => ddr_dqs_to_and_from_the_ddr_sdram_0,
      ddr_ras_n => internal_ddr_ras_n_from_the_ddr_sdram_0,
      ddr_we_n => internal_ddr_we_n_from_the_ddr_sdram_0,
      local_rdata => ddr_sdram_0_s1_readdata,
      local_rdata_valid => ddr_sdram_0_s1_readdatavalid,
      local_ready => ddr_sdram_0_s1_waitrequest_n,
      stratix_dll_control => internal_stratix_dll_control_from_the_ddr_sdram_0,
      clk => internal_pll_c0_out,
      dqs_delay_ctrl => dqs_delay_ctrl_to_the_ddr_sdram_0,
      dqsupdate => dqsupdate_to_the_ddr_sdram_0,
      local_addr => ddr_sdram_0_s1_address,
      local_be => ddr_sdram_0_s1_byteenable,
      local_read_req => ddr_sdram_0_s1_read,
      local_wdata => ddr_sdram_0_s1_writedata,
      local_write_req => ddr_sdram_0_s1_write,
      reset_n => ddr_sdram_0_s1_reset_n,
      write_clk => write_clk_to_the_ddr_sdram_0
    );


  --the_descriptor_memory_s1, which is an e_instance
  the_descriptor_memory_s1 : descriptor_memory_s1_arbitrator
    port map(
      cpu_data_master_granted_descriptor_memory_s1 => cpu_data_master_granted_descriptor_memory_s1,
      cpu_data_master_qualified_request_descriptor_memory_s1 => cpu_data_master_qualified_request_descriptor_memory_s1,
      cpu_data_master_read_data_valid_descriptor_memory_s1 => cpu_data_master_read_data_valid_descriptor_memory_s1,
      cpu_data_master_requests_descriptor_memory_s1 => cpu_data_master_requests_descriptor_memory_s1,
      d1_descriptor_memory_s1_end_xfer => d1_descriptor_memory_s1_end_xfer,
      descriptor_memory_s1_address => descriptor_memory_s1_address,
      descriptor_memory_s1_byteenable => descriptor_memory_s1_byteenable,
      descriptor_memory_s1_chipselect => descriptor_memory_s1_chipselect,
      descriptor_memory_s1_clken => descriptor_memory_s1_clken,
      descriptor_memory_s1_readdata_from_sa => descriptor_memory_s1_readdata_from_sa,
      descriptor_memory_s1_write => descriptor_memory_s1_write,
      descriptor_memory_s1_writedata => descriptor_memory_s1_writedata,
      sgdma_rx_descriptor_read_granted_descriptor_memory_s1 => sgdma_rx_descriptor_read_granted_descriptor_memory_s1,
      sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 => sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1,
      sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1 => sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1,
      sgdma_rx_descriptor_read_requests_descriptor_memory_s1 => sgdma_rx_descriptor_read_requests_descriptor_memory_s1,
      sgdma_rx_descriptor_write_granted_descriptor_memory_s1 => sgdma_rx_descriptor_write_granted_descriptor_memory_s1,
      sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 => sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1,
      sgdma_rx_descriptor_write_requests_descriptor_memory_s1 => sgdma_rx_descriptor_write_requests_descriptor_memory_s1,
      sgdma_tx_descriptor_read_granted_descriptor_memory_s1 => sgdma_tx_descriptor_read_granted_descriptor_memory_s1,
      sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 => sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1,
      sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1 => sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1,
      sgdma_tx_descriptor_read_requests_descriptor_memory_s1 => sgdma_tx_descriptor_read_requests_descriptor_memory_s1,
      sgdma_tx_descriptor_write_granted_descriptor_memory_s1 => sgdma_tx_descriptor_write_granted_descriptor_memory_s1,
      sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 => sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1,
      sgdma_tx_descriptor_write_requests_descriptor_memory_s1 => sgdma_tx_descriptor_write_requests_descriptor_memory_s1,
      clk => internal_pll_c0_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      descriptor_memory_s1_readdata => descriptor_memory_s1_readdata,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_descriptor_read_address_to_slave => sgdma_rx_descriptor_read_address_to_slave,
      sgdma_rx_descriptor_read_latency_counter => sgdma_rx_descriptor_read_latency_counter,
      sgdma_rx_descriptor_read_read => sgdma_rx_descriptor_read_read,
      sgdma_rx_descriptor_write_address_to_slave => sgdma_rx_descriptor_write_address_to_slave,
      sgdma_rx_descriptor_write_write => sgdma_rx_descriptor_write_write,
      sgdma_rx_descriptor_write_writedata => sgdma_rx_descriptor_write_writedata,
      sgdma_tx_descriptor_read_address_to_slave => sgdma_tx_descriptor_read_address_to_slave,
      sgdma_tx_descriptor_read_latency_counter => sgdma_tx_descriptor_read_latency_counter,
      sgdma_tx_descriptor_read_read => sgdma_tx_descriptor_read_read,
      sgdma_tx_descriptor_write_address_to_slave => sgdma_tx_descriptor_write_address_to_slave,
      sgdma_tx_descriptor_write_write => sgdma_tx_descriptor_write_write,
      sgdma_tx_descriptor_write_writedata => sgdma_tx_descriptor_write_writedata
    );


  --the_descriptor_memory, which is an e_ptf_instance
  the_descriptor_memory : descriptor_memory
    port map(
      readdata => descriptor_memory_s1_readdata,
      address => descriptor_memory_s1_address,
      byteenable => descriptor_memory_s1_byteenable,
      chipselect => descriptor_memory_s1_chipselect,
      clk => internal_pll_c0_out,
      clken => descriptor_memory_s1_clken,
      write => descriptor_memory_s1_write,
      writedata => descriptor_memory_s1_writedata
    );


  --the_ext_flash_enet_bus_avalon_slave, which is an e_instance
  the_ext_flash_enet_bus_avalon_slave : ext_flash_enet_bus_avalon_slave_arbitrator
    port map(
      d1_ext_flash_enet_bus_avalon_slave_end_xfer => d1_ext_flash_enet_bus_avalon_slave_end_xfer,
      ext_flash_enet_bus_address => internal_ext_flash_enet_bus_address,
      ext_flash_enet_bus_data => ext_flash_enet_bus_data,
      ext_flash_s1_wait_counter_eq_0 => ext_flash_s1_wait_counter_eq_0,
      incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0 => incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0,
      pipeline_bridge_m1_byteenable_ext_flash_s1 => pipeline_bridge_m1_byteenable_ext_flash_s1,
      pipeline_bridge_m1_granted_ext_flash_s1 => pipeline_bridge_m1_granted_ext_flash_s1,
      pipeline_bridge_m1_qualified_request_ext_flash_s1 => pipeline_bridge_m1_qualified_request_ext_flash_s1,
      pipeline_bridge_m1_read_data_valid_ext_flash_s1 => pipeline_bridge_m1_read_data_valid_ext_flash_s1,
      pipeline_bridge_m1_requests_ext_flash_s1 => pipeline_bridge_m1_requests_ext_flash_s1,
      read_n_to_the_ext_flash => internal_read_n_to_the_ext_flash,
      select_n_to_the_ext_flash => internal_select_n_to_the_ext_flash,
      write_n_to_the_ext_flash => internal_write_n_to_the_ext_flash,
      clk => internal_pll_c0_out,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_byteenable => pipeline_bridge_m1_byteenable,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_dbs_address => pipeline_bridge_m1_dbs_address,
      pipeline_bridge_m1_dbs_write_8 => pipeline_bridge_m1_dbs_write_8,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      reset_n => pll_c0_out_reset_n
    );


  --the_ext_ssram_bus_avalon_slave, which is an e_instance
  the_ext_ssram_bus_avalon_slave : ext_ssram_bus_avalon_slave_arbitrator
    port map(
      adsc_n_to_the_ext_ssram => internal_adsc_n_to_the_ext_ssram,
      bw_n_to_the_ext_ssram => internal_bw_n_to_the_ext_ssram,
      bwe_n_to_the_ext_ssram => internal_bwe_n_to_the_ext_ssram,
      chipenable1_n_to_the_ext_ssram => internal_chipenable1_n_to_the_ext_ssram,
      cpu_data_master_granted_ext_ssram_s1 => cpu_data_master_granted_ext_ssram_s1,
      cpu_data_master_qualified_request_ext_ssram_s1 => cpu_data_master_qualified_request_ext_ssram_s1,
      cpu_data_master_read_data_valid_ext_ssram_s1 => cpu_data_master_read_data_valid_ext_ssram_s1,
      cpu_data_master_requests_ext_ssram_s1 => cpu_data_master_requests_ext_ssram_s1,
      cpu_instruction_master_granted_ext_ssram_s1 => cpu_instruction_master_granted_ext_ssram_s1,
      cpu_instruction_master_qualified_request_ext_ssram_s1 => cpu_instruction_master_qualified_request_ext_ssram_s1,
      cpu_instruction_master_read_data_valid_ext_ssram_s1 => cpu_instruction_master_read_data_valid_ext_ssram_s1,
      cpu_instruction_master_requests_ext_ssram_s1 => cpu_instruction_master_requests_ext_ssram_s1,
      d1_ext_ssram_bus_avalon_slave_end_xfer => d1_ext_ssram_bus_avalon_slave_end_xfer,
      ext_ssram_bus_address => internal_ext_ssram_bus_address,
      ext_ssram_bus_data => ext_ssram_bus_data,
      incoming_ext_ssram_bus_data => incoming_ext_ssram_bus_data,
      outputenable_n_to_the_ext_ssram => internal_outputenable_n_to_the_ext_ssram,
      sgdma_rx_m_write_granted_ext_ssram_s1 => sgdma_rx_m_write_granted_ext_ssram_s1,
      sgdma_rx_m_write_qualified_request_ext_ssram_s1 => sgdma_rx_m_write_qualified_request_ext_ssram_s1,
      sgdma_rx_m_write_requests_ext_ssram_s1 => sgdma_rx_m_write_requests_ext_ssram_s1,
      sgdma_tx_m_read_granted_ext_ssram_s1 => sgdma_tx_m_read_granted_ext_ssram_s1,
      sgdma_tx_m_read_qualified_request_ext_ssram_s1 => sgdma_tx_m_read_qualified_request_ext_ssram_s1,
      sgdma_tx_m_read_read_data_valid_ext_ssram_s1 => sgdma_tx_m_read_read_data_valid_ext_ssram_s1,
      sgdma_tx_m_read_requests_ext_ssram_s1 => sgdma_tx_m_read_requests_ext_ssram_s1,
      clk => internal_pll_c0_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_m_write_address_to_slave => sgdma_rx_m_write_address_to_slave,
      sgdma_rx_m_write_byteenable => sgdma_rx_m_write_byteenable,
      sgdma_rx_m_write_write => sgdma_rx_m_write_write,
      sgdma_rx_m_write_writedata => sgdma_rx_m_write_writedata,
      sgdma_tx_m_read_address_to_slave => sgdma_tx_m_read_address_to_slave,
      sgdma_tx_m_read_latency_counter => sgdma_tx_m_read_latency_counter,
      sgdma_tx_m_read_read => sgdma_tx_m_read_read,
      sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register => sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register
    );


  --the_high_res_timer_s1, which is an e_instance
  the_high_res_timer_s1 : high_res_timer_s1_arbitrator
    port map(
      d1_high_res_timer_s1_end_xfer => d1_high_res_timer_s1_end_xfer,
      high_res_timer_s1_address => high_res_timer_s1_address,
      high_res_timer_s1_chipselect => high_res_timer_s1_chipselect,
      high_res_timer_s1_irq_from_sa => high_res_timer_s1_irq_from_sa,
      high_res_timer_s1_readdata_from_sa => high_res_timer_s1_readdata_from_sa,
      high_res_timer_s1_reset_n => high_res_timer_s1_reset_n,
      high_res_timer_s1_write_n => high_res_timer_s1_write_n,
      high_res_timer_s1_writedata => high_res_timer_s1_writedata,
      pipeline_bridge_m1_granted_high_res_timer_s1 => pipeline_bridge_m1_granted_high_res_timer_s1,
      pipeline_bridge_m1_qualified_request_high_res_timer_s1 => pipeline_bridge_m1_qualified_request_high_res_timer_s1,
      pipeline_bridge_m1_read_data_valid_high_res_timer_s1 => pipeline_bridge_m1_read_data_valid_high_res_timer_s1,
      pipeline_bridge_m1_requests_high_res_timer_s1 => pipeline_bridge_m1_requests_high_res_timer_s1,
      clk => internal_pll_c0_out,
      high_res_timer_s1_irq => high_res_timer_s1_irq,
      high_res_timer_s1_readdata => high_res_timer_s1_readdata,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n
    );


  --the_high_res_timer, which is an e_ptf_instance
  the_high_res_timer : high_res_timer
    port map(
      irq => high_res_timer_s1_irq,
      readdata => high_res_timer_s1_readdata,
      address => high_res_timer_s1_address,
      chipselect => high_res_timer_s1_chipselect,
      clk => internal_pll_c0_out,
      reset_n => high_res_timer_s1_reset_n,
      write_n => high_res_timer_s1_write_n,
      writedata => high_res_timer_s1_writedata
    );


  --the_interrupt_vector_interrupt_vector, which is an e_instance
  the_interrupt_vector_interrupt_vector : interrupt_vector_interrupt_vector_arbitrator
    port map(
      interrupt_vector_interrupt_vector_estatus => interrupt_vector_interrupt_vector_estatus,
      interrupt_vector_interrupt_vector_ipending => interrupt_vector_interrupt_vector_ipending,
      interrupt_vector_interrupt_vector_result_from_sa => interrupt_vector_interrupt_vector_result_from_sa,
      clk => internal_pll_c0_out,
      cpu_custom_instruction_master_combo_estatus => cpu_custom_instruction_master_combo_estatus,
      cpu_custom_instruction_master_combo_ipending => cpu_custom_instruction_master_combo_ipending,
      interrupt_vector_interrupt_vector_result => interrupt_vector_interrupt_vector_result,
      interrupt_vector_interrupt_vector_select => interrupt_vector_interrupt_vector_select,
      reset_n => pll_c0_out_reset_n
    );


  --the_interrupt_vector, which is an e_ptf_instance
  the_interrupt_vector : interrupt_vector
    port map(
      result => interrupt_vector_interrupt_vector_result,
      estatus => interrupt_vector_interrupt_vector_estatus,
      ipending => interrupt_vector_interrupt_vector_ipending
    );


  --the_jtag_uart_avalon_jtag_slave, which is an e_instance
  the_jtag_uart_avalon_jtag_slave : jtag_uart_avalon_jtag_slave_arbitrator
    port map(
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      jtag_uart_avalon_jtag_slave_address => jtag_uart_avalon_jtag_slave_address,
      jtag_uart_avalon_jtag_slave_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      jtag_uart_avalon_jtag_slave_dataavailable_from_sa => jtag_uart_avalon_jtag_slave_dataavailable_from_sa,
      jtag_uart_avalon_jtag_slave_irq_from_sa => jtag_uart_avalon_jtag_slave_irq_from_sa,
      jtag_uart_avalon_jtag_slave_read_n => jtag_uart_avalon_jtag_slave_read_n,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_readyfordata_from_sa => jtag_uart_avalon_jtag_slave_readyfordata_from_sa,
      jtag_uart_avalon_jtag_slave_reset_n => jtag_uart_avalon_jtag_slave_reset_n,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      jtag_uart_avalon_jtag_slave_write_n => jtag_uart_avalon_jtag_slave_write_n,
      jtag_uart_avalon_jtag_slave_writedata => jtag_uart_avalon_jtag_slave_writedata,
      pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave => pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave,
      pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave => pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave,
      pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave => pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
      pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave => pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave,
      clk => internal_pll_c0_out,
      jtag_uart_avalon_jtag_slave_dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      jtag_uart_avalon_jtag_slave_irq => jtag_uart_avalon_jtag_slave_irq,
      jtag_uart_avalon_jtag_slave_readdata => jtag_uart_avalon_jtag_slave_readdata,
      jtag_uart_avalon_jtag_slave_readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      jtag_uart_avalon_jtag_slave_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n
    );


  --the_jtag_uart, which is an e_ptf_instance
  the_jtag_uart : jtag_uart
    port map(
      av_irq => jtag_uart_avalon_jtag_slave_irq,
      av_readdata => jtag_uart_avalon_jtag_slave_readdata,
      av_waitrequest => jtag_uart_avalon_jtag_slave_waitrequest,
      dataavailable => jtag_uart_avalon_jtag_slave_dataavailable,
      readyfordata => jtag_uart_avalon_jtag_slave_readyfordata,
      av_address => jtag_uart_avalon_jtag_slave_address,
      av_chipselect => jtag_uart_avalon_jtag_slave_chipselect,
      av_read_n => jtag_uart_avalon_jtag_slave_read_n,
      av_write_n => jtag_uart_avalon_jtag_slave_write_n,
      av_writedata => jtag_uart_avalon_jtag_slave_writedata,
      clk => internal_pll_c0_out,
      rst_n => jtag_uart_avalon_jtag_slave_reset_n
    );


  --the_lcd_display_control_slave, which is an e_instance
  the_lcd_display_control_slave : lcd_display_control_slave_arbitrator
    port map(
      d1_lcd_display_control_slave_end_xfer => d1_lcd_display_control_slave_end_xfer,
      lcd_display_control_slave_address => lcd_display_control_slave_address,
      lcd_display_control_slave_begintransfer => lcd_display_control_slave_begintransfer,
      lcd_display_control_slave_read => lcd_display_control_slave_read,
      lcd_display_control_slave_readdata_from_sa => lcd_display_control_slave_readdata_from_sa,
      lcd_display_control_slave_wait_counter_eq_0 => lcd_display_control_slave_wait_counter_eq_0,
      lcd_display_control_slave_write => lcd_display_control_slave_write,
      lcd_display_control_slave_writedata => lcd_display_control_slave_writedata,
      pipeline_bridge_m1_granted_lcd_display_control_slave => pipeline_bridge_m1_granted_lcd_display_control_slave,
      pipeline_bridge_m1_qualified_request_lcd_display_control_slave => pipeline_bridge_m1_qualified_request_lcd_display_control_slave,
      pipeline_bridge_m1_read_data_valid_lcd_display_control_slave => pipeline_bridge_m1_read_data_valid_lcd_display_control_slave,
      pipeline_bridge_m1_requests_lcd_display_control_slave => pipeline_bridge_m1_requests_lcd_display_control_slave,
      clk => internal_pll_c0_out,
      lcd_display_control_slave_readdata => lcd_display_control_slave_readdata,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_byteenable => pipeline_bridge_m1_byteenable,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n
    );


  --the_lcd_display, which is an e_ptf_instance
  the_lcd_display : lcd_display
    port map(
      LCD_E => internal_LCD_E_from_the_lcd_display,
      LCD_RS => internal_LCD_RS_from_the_lcd_display,
      LCD_RW => internal_LCD_RW_from_the_lcd_display,
      LCD_data => LCD_data_to_and_from_the_lcd_display,
      readdata => lcd_display_control_slave_readdata,
      address => lcd_display_control_slave_address,
      begintransfer => lcd_display_control_slave_begintransfer,
      read => lcd_display_control_slave_read,
      write => lcd_display_control_slave_write,
      writedata => lcd_display_control_slave_writedata
    );


  --the_led_pio_s1, which is an e_instance
  the_led_pio_s1 : led_pio_s1_arbitrator
    port map(
      d1_led_pio_s1_end_xfer => d1_led_pio_s1_end_xfer,
      led_pio_s1_address => led_pio_s1_address,
      led_pio_s1_chipselect => led_pio_s1_chipselect,
      led_pio_s1_readdata_from_sa => led_pio_s1_readdata_from_sa,
      led_pio_s1_reset_n => led_pio_s1_reset_n,
      led_pio_s1_write_n => led_pio_s1_write_n,
      led_pio_s1_writedata => led_pio_s1_writedata,
      pipeline_bridge_m1_granted_led_pio_s1 => pipeline_bridge_m1_granted_led_pio_s1,
      pipeline_bridge_m1_qualified_request_led_pio_s1 => pipeline_bridge_m1_qualified_request_led_pio_s1,
      pipeline_bridge_m1_read_data_valid_led_pio_s1 => pipeline_bridge_m1_read_data_valid_led_pio_s1,
      pipeline_bridge_m1_requests_led_pio_s1 => pipeline_bridge_m1_requests_led_pio_s1,
      clk => internal_pll_c0_out,
      led_pio_s1_readdata => led_pio_s1_readdata,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_byteenable => pipeline_bridge_m1_byteenable,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n
    );


  --the_led_pio, which is an e_ptf_instance
  the_led_pio : led_pio
    port map(
      out_port => internal_out_port_from_the_led_pio,
      readdata => led_pio_s1_readdata,
      address => led_pio_s1_address,
      chipselect => led_pio_s1_chipselect,
      clk => internal_pll_c0_out,
      reset_n => led_pio_s1_reset_n,
      write_n => led_pio_s1_write_n,
      writedata => led_pio_s1_writedata
    );


  --the_packet_memory_s1, which is an e_instance
  the_packet_memory_s1 : packet_memory_s1_arbitrator
    port map(
      cpu_data_master_granted_packet_memory_s1 => cpu_data_master_granted_packet_memory_s1,
      cpu_data_master_qualified_request_packet_memory_s1 => cpu_data_master_qualified_request_packet_memory_s1,
      cpu_data_master_read_data_valid_packet_memory_s1 => cpu_data_master_read_data_valid_packet_memory_s1,
      cpu_data_master_requests_packet_memory_s1 => cpu_data_master_requests_packet_memory_s1,
      d1_packet_memory_s1_end_xfer => d1_packet_memory_s1_end_xfer,
      packet_memory_s1_address => packet_memory_s1_address,
      packet_memory_s1_byteenable => packet_memory_s1_byteenable,
      packet_memory_s1_chipselect => packet_memory_s1_chipselect,
      packet_memory_s1_clken => packet_memory_s1_clken,
      packet_memory_s1_readdata_from_sa => packet_memory_s1_readdata_from_sa,
      packet_memory_s1_write => packet_memory_s1_write,
      packet_memory_s1_writedata => packet_memory_s1_writedata,
      clk => internal_pll_c0_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      packet_memory_s1_readdata => packet_memory_s1_readdata,
      reset_n => pll_c0_out_reset_n
    );


  --the_packet_memory_s2, which is an e_instance
  the_packet_memory_s2 : packet_memory_s2_arbitrator
    port map(
      d1_packet_memory_s2_end_xfer => d1_packet_memory_s2_end_xfer,
      packet_memory_s2_address => packet_memory_s2_address,
      packet_memory_s2_byteenable => packet_memory_s2_byteenable,
      packet_memory_s2_chipselect => packet_memory_s2_chipselect,
      packet_memory_s2_clken => packet_memory_s2_clken,
      packet_memory_s2_readdata_from_sa => packet_memory_s2_readdata_from_sa,
      packet_memory_s2_write => packet_memory_s2_write,
      packet_memory_s2_writedata => packet_memory_s2_writedata,
      sgdma_rx_m_write_granted_packet_memory_s2 => sgdma_rx_m_write_granted_packet_memory_s2,
      sgdma_rx_m_write_qualified_request_packet_memory_s2 => sgdma_rx_m_write_qualified_request_packet_memory_s2,
      sgdma_rx_m_write_requests_packet_memory_s2 => sgdma_rx_m_write_requests_packet_memory_s2,
      sgdma_tx_m_read_granted_packet_memory_s2 => sgdma_tx_m_read_granted_packet_memory_s2,
      sgdma_tx_m_read_qualified_request_packet_memory_s2 => sgdma_tx_m_read_qualified_request_packet_memory_s2,
      sgdma_tx_m_read_read_data_valid_packet_memory_s2 => sgdma_tx_m_read_read_data_valid_packet_memory_s2,
      sgdma_tx_m_read_requests_packet_memory_s2 => sgdma_tx_m_read_requests_packet_memory_s2,
      clk => internal_pll_c0_out,
      packet_memory_s2_readdata => packet_memory_s2_readdata,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_m_write_address_to_slave => sgdma_rx_m_write_address_to_slave,
      sgdma_rx_m_write_byteenable => sgdma_rx_m_write_byteenable,
      sgdma_rx_m_write_write => sgdma_rx_m_write_write,
      sgdma_rx_m_write_writedata => sgdma_rx_m_write_writedata,
      sgdma_tx_m_read_address_to_slave => sgdma_tx_m_read_address_to_slave,
      sgdma_tx_m_read_latency_counter => sgdma_tx_m_read_latency_counter,
      sgdma_tx_m_read_read => sgdma_tx_m_read_read,
      sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register => sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register
    );


  --the_packet_memory, which is an e_ptf_instance
  the_packet_memory : packet_memory
    port map(
      readdata => packet_memory_s1_readdata,
      readdata2 => packet_memory_s2_readdata,
      address => packet_memory_s1_address,
      address2 => packet_memory_s2_address,
      byteenable => packet_memory_s1_byteenable,
      byteenable2 => packet_memory_s2_byteenable,
      chipselect => packet_memory_s1_chipselect,
      chipselect2 => packet_memory_s2_chipselect,
      clk => internal_pll_c0_out,
      clk2 => internal_pll_c0_out,
      clken => packet_memory_s1_clken,
      clken2 => packet_memory_s2_clken,
      write => packet_memory_s1_write,
      write2 => packet_memory_s2_write,
      writedata => packet_memory_s1_writedata,
      writedata2 => packet_memory_s2_writedata
    );


  --the_pipeline_bridge_s1, which is an e_instance
  the_pipeline_bridge_s1 : pipeline_bridge_s1_arbitrator
    port map(
      cpu_data_master_granted_pipeline_bridge_s1 => cpu_data_master_granted_pipeline_bridge_s1,
      cpu_data_master_qualified_request_pipeline_bridge_s1 => cpu_data_master_qualified_request_pipeline_bridge_s1,
      cpu_data_master_read_data_valid_pipeline_bridge_s1 => cpu_data_master_read_data_valid_pipeline_bridge_s1,
      cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register,
      cpu_data_master_requests_pipeline_bridge_s1 => cpu_data_master_requests_pipeline_bridge_s1,
      cpu_instruction_master_granted_pipeline_bridge_s1 => cpu_instruction_master_granted_pipeline_bridge_s1,
      cpu_instruction_master_qualified_request_pipeline_bridge_s1 => cpu_instruction_master_qualified_request_pipeline_bridge_s1,
      cpu_instruction_master_read_data_valid_pipeline_bridge_s1 => cpu_instruction_master_read_data_valid_pipeline_bridge_s1,
      cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_instruction_master_read_data_valid_pipeline_bridge_s1_shift_register,
      cpu_instruction_master_requests_pipeline_bridge_s1 => cpu_instruction_master_requests_pipeline_bridge_s1,
      d1_pipeline_bridge_s1_end_xfer => d1_pipeline_bridge_s1_end_xfer,
      pipeline_bridge_s1_address => pipeline_bridge_s1_address,
      pipeline_bridge_s1_arbiterlock => pipeline_bridge_s1_arbiterlock,
      pipeline_bridge_s1_arbiterlock2 => pipeline_bridge_s1_arbiterlock2,
      pipeline_bridge_s1_burstcount => pipeline_bridge_s1_burstcount,
      pipeline_bridge_s1_byteenable => pipeline_bridge_s1_byteenable,
      pipeline_bridge_s1_chipselect => pipeline_bridge_s1_chipselect,
      pipeline_bridge_s1_debugaccess => pipeline_bridge_s1_debugaccess,
      pipeline_bridge_s1_endofpacket_from_sa => pipeline_bridge_s1_endofpacket_from_sa,
      pipeline_bridge_s1_nativeaddress => pipeline_bridge_s1_nativeaddress,
      pipeline_bridge_s1_read => pipeline_bridge_s1_read,
      pipeline_bridge_s1_readdata_from_sa => pipeline_bridge_s1_readdata_from_sa,
      pipeline_bridge_s1_reset_n => pipeline_bridge_s1_reset_n,
      pipeline_bridge_s1_waitrequest_from_sa => pipeline_bridge_s1_waitrequest_from_sa,
      pipeline_bridge_s1_write => pipeline_bridge_s1_write,
      pipeline_bridge_s1_writedata => pipeline_bridge_s1_writedata,
      clk => internal_pll_c0_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_byteenable => cpu_data_master_byteenable,
      cpu_data_master_debugaccess => cpu_data_master_debugaccess,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      cpu_instruction_master_address_to_slave => cpu_instruction_master_address_to_slave,
      cpu_instruction_master_latency_counter => cpu_instruction_master_latency_counter,
      cpu_instruction_master_read => cpu_instruction_master_read,
      cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_instruction_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      pipeline_bridge_s1_endofpacket => pipeline_bridge_s1_endofpacket,
      pipeline_bridge_s1_readdata => pipeline_bridge_s1_readdata,
      pipeline_bridge_s1_readdatavalid => pipeline_bridge_s1_readdatavalid,
      pipeline_bridge_s1_waitrequest => pipeline_bridge_s1_waitrequest,
      reset_n => pll_c0_out_reset_n
    );


  --the_pipeline_bridge_m1, which is an e_instance
  the_pipeline_bridge_m1 : pipeline_bridge_m1_arbitrator
    port map(
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_dbs_address => pipeline_bridge_m1_dbs_address,
      pipeline_bridge_m1_dbs_write_8 => pipeline_bridge_m1_dbs_write_8,
      pipeline_bridge_m1_endofpacket => pipeline_bridge_m1_endofpacket,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_readdata => pipeline_bridge_m1_readdata,
      pipeline_bridge_m1_readdatavalid => pipeline_bridge_m1_readdatavalid,
      pipeline_bridge_m1_waitrequest => pipeline_bridge_m1_waitrequest,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_endofpacket_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_readdata_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_waitrequest_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_endofpacket_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_readdata_from_sa,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_waitrequest_from_sa,
      button_pio_s1_readdata_from_sa => button_pio_s1_readdata_from_sa,
      clk => internal_pll_c0_out,
      cpu_jtag_debug_module_readdata_from_sa => cpu_jtag_debug_module_readdata_from_sa,
      d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer => d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in_end_xfer,
      d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer => d1_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in_end_xfer,
      d1_button_pio_s1_end_xfer => d1_button_pio_s1_end_xfer,
      d1_cpu_jtag_debug_module_end_xfer => d1_cpu_jtag_debug_module_end_xfer,
      d1_ext_flash_enet_bus_avalon_slave_end_xfer => d1_ext_flash_enet_bus_avalon_slave_end_xfer,
      d1_high_res_timer_s1_end_xfer => d1_high_res_timer_s1_end_xfer,
      d1_jtag_uart_avalon_jtag_slave_end_xfer => d1_jtag_uart_avalon_jtag_slave_end_xfer,
      d1_lcd_display_control_slave_end_xfer => d1_lcd_display_control_slave_end_xfer,
      d1_led_pio_s1_end_xfer => d1_led_pio_s1_end_xfer,
      d1_reconfig_request_pio_s1_end_xfer => d1_reconfig_request_pio_s1_end_xfer,
      d1_seven_seg_pio_s1_end_xfer => d1_seven_seg_pio_s1_end_xfer,
      d1_sgdma_rx_csr_end_xfer => d1_sgdma_rx_csr_end_xfer,
      d1_sgdma_tx_csr_end_xfer => d1_sgdma_tx_csr_end_xfer,
      d1_sys_clk_timer_s1_end_xfer => d1_sys_clk_timer_s1_end_xfer,
      d1_uart1_s1_end_xfer => d1_uart1_s1_end_xfer,
      ext_flash_s1_wait_counter_eq_0 => ext_flash_s1_wait_counter_eq_0,
      high_res_timer_s1_readdata_from_sa => high_res_timer_s1_readdata_from_sa,
      incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0 => incoming_ext_flash_enet_bus_data_with_Xs_converted_to_0,
      jtag_uart_avalon_jtag_slave_readdata_from_sa => jtag_uart_avalon_jtag_slave_readdata_from_sa,
      jtag_uart_avalon_jtag_slave_waitrequest_from_sa => jtag_uart_avalon_jtag_slave_waitrequest_from_sa,
      lcd_display_control_slave_readdata_from_sa => lcd_display_control_slave_readdata_from_sa,
      lcd_display_control_slave_wait_counter_eq_0 => lcd_display_control_slave_wait_counter_eq_0,
      led_pio_s1_readdata_from_sa => led_pio_s1_readdata_from_sa,
      pipeline_bridge_m1_address => pipeline_bridge_m1_address,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_byteenable => pipeline_bridge_m1_byteenable,
      pipeline_bridge_m1_byteenable_ext_flash_s1 => pipeline_bridge_m1_byteenable_ext_flash_s1,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in => pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in,
      pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in => pipeline_bridge_m1_granted_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in,
      pipeline_bridge_m1_granted_button_pio_s1 => pipeline_bridge_m1_granted_button_pio_s1,
      pipeline_bridge_m1_granted_cpu_jtag_debug_module => pipeline_bridge_m1_granted_cpu_jtag_debug_module,
      pipeline_bridge_m1_granted_ext_flash_s1 => pipeline_bridge_m1_granted_ext_flash_s1,
      pipeline_bridge_m1_granted_high_res_timer_s1 => pipeline_bridge_m1_granted_high_res_timer_s1,
      pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave => pipeline_bridge_m1_granted_jtag_uart_avalon_jtag_slave,
      pipeline_bridge_m1_granted_lcd_display_control_slave => pipeline_bridge_m1_granted_lcd_display_control_slave,
      pipeline_bridge_m1_granted_led_pio_s1 => pipeline_bridge_m1_granted_led_pio_s1,
      pipeline_bridge_m1_granted_reconfig_request_pio_s1 => pipeline_bridge_m1_granted_reconfig_request_pio_s1,
      pipeline_bridge_m1_granted_seven_seg_pio_s1 => pipeline_bridge_m1_granted_seven_seg_pio_s1,
      pipeline_bridge_m1_granted_sgdma_rx_csr => pipeline_bridge_m1_granted_sgdma_rx_csr,
      pipeline_bridge_m1_granted_sgdma_tx_csr => pipeline_bridge_m1_granted_sgdma_tx_csr,
      pipeline_bridge_m1_granted_sys_clk_timer_s1 => pipeline_bridge_m1_granted_sys_clk_timer_s1,
      pipeline_bridge_m1_granted_uart1_s1 => pipeline_bridge_m1_granted_uart1_s1,
      pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in => pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in,
      pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in => pipeline_bridge_m1_qualified_request_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in,
      pipeline_bridge_m1_qualified_request_button_pio_s1 => pipeline_bridge_m1_qualified_request_button_pio_s1,
      pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module => pipeline_bridge_m1_qualified_request_cpu_jtag_debug_module,
      pipeline_bridge_m1_qualified_request_ext_flash_s1 => pipeline_bridge_m1_qualified_request_ext_flash_s1,
      pipeline_bridge_m1_qualified_request_high_res_timer_s1 => pipeline_bridge_m1_qualified_request_high_res_timer_s1,
      pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave => pipeline_bridge_m1_qualified_request_jtag_uart_avalon_jtag_slave,
      pipeline_bridge_m1_qualified_request_lcd_display_control_slave => pipeline_bridge_m1_qualified_request_lcd_display_control_slave,
      pipeline_bridge_m1_qualified_request_led_pio_s1 => pipeline_bridge_m1_qualified_request_led_pio_s1,
      pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 => pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1,
      pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 => pipeline_bridge_m1_qualified_request_seven_seg_pio_s1,
      pipeline_bridge_m1_qualified_request_sgdma_rx_csr => pipeline_bridge_m1_qualified_request_sgdma_rx_csr,
      pipeline_bridge_m1_qualified_request_sgdma_tx_csr => pipeline_bridge_m1_qualified_request_sgdma_tx_csr,
      pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 => pipeline_bridge_m1_qualified_request_sys_clk_timer_s1,
      pipeline_bridge_m1_qualified_request_uart1_s1 => pipeline_bridge_m1_qualified_request_uart1_s1,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in => pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in,
      pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in => pipeline_bridge_m1_read_data_valid_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in,
      pipeline_bridge_m1_read_data_valid_button_pio_s1 => pipeline_bridge_m1_read_data_valid_button_pio_s1,
      pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module => pipeline_bridge_m1_read_data_valid_cpu_jtag_debug_module,
      pipeline_bridge_m1_read_data_valid_ext_flash_s1 => pipeline_bridge_m1_read_data_valid_ext_flash_s1,
      pipeline_bridge_m1_read_data_valid_high_res_timer_s1 => pipeline_bridge_m1_read_data_valid_high_res_timer_s1,
      pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave => pipeline_bridge_m1_read_data_valid_jtag_uart_avalon_jtag_slave,
      pipeline_bridge_m1_read_data_valid_lcd_display_control_slave => pipeline_bridge_m1_read_data_valid_lcd_display_control_slave,
      pipeline_bridge_m1_read_data_valid_led_pio_s1 => pipeline_bridge_m1_read_data_valid_led_pio_s1,
      pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1 => pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1,
      pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1 => pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1,
      pipeline_bridge_m1_read_data_valid_sgdma_rx_csr => pipeline_bridge_m1_read_data_valid_sgdma_rx_csr,
      pipeline_bridge_m1_read_data_valid_sgdma_tx_csr => pipeline_bridge_m1_read_data_valid_sgdma_tx_csr,
      pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1 => pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1,
      pipeline_bridge_m1_read_data_valid_uart1_s1 => pipeline_bridge_m1_read_data_valid_uart1_s1,
      pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in => pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_in,
      pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in => pipeline_bridge_m1_requests_NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_in,
      pipeline_bridge_m1_requests_button_pio_s1 => pipeline_bridge_m1_requests_button_pio_s1,
      pipeline_bridge_m1_requests_cpu_jtag_debug_module => pipeline_bridge_m1_requests_cpu_jtag_debug_module,
      pipeline_bridge_m1_requests_ext_flash_s1 => pipeline_bridge_m1_requests_ext_flash_s1,
      pipeline_bridge_m1_requests_high_res_timer_s1 => pipeline_bridge_m1_requests_high_res_timer_s1,
      pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave => pipeline_bridge_m1_requests_jtag_uart_avalon_jtag_slave,
      pipeline_bridge_m1_requests_lcd_display_control_slave => pipeline_bridge_m1_requests_lcd_display_control_slave,
      pipeline_bridge_m1_requests_led_pio_s1 => pipeline_bridge_m1_requests_led_pio_s1,
      pipeline_bridge_m1_requests_reconfig_request_pio_s1 => pipeline_bridge_m1_requests_reconfig_request_pio_s1,
      pipeline_bridge_m1_requests_seven_seg_pio_s1 => pipeline_bridge_m1_requests_seven_seg_pio_s1,
      pipeline_bridge_m1_requests_sgdma_rx_csr => pipeline_bridge_m1_requests_sgdma_rx_csr,
      pipeline_bridge_m1_requests_sgdma_tx_csr => pipeline_bridge_m1_requests_sgdma_tx_csr,
      pipeline_bridge_m1_requests_sys_clk_timer_s1 => pipeline_bridge_m1_requests_sys_clk_timer_s1,
      pipeline_bridge_m1_requests_uart1_s1 => pipeline_bridge_m1_requests_uart1_s1,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reconfig_request_pio_s1_readdata_from_sa => reconfig_request_pio_s1_readdata_from_sa,
      reset_n => pll_c0_out_reset_n,
      seven_seg_pio_s1_readdata_from_sa => seven_seg_pio_s1_readdata_from_sa,
      sgdma_rx_csr_readdata_from_sa => sgdma_rx_csr_readdata_from_sa,
      sgdma_tx_csr_readdata_from_sa => sgdma_tx_csr_readdata_from_sa,
      sys_clk_timer_s1_readdata_from_sa => sys_clk_timer_s1_readdata_from_sa,
      uart1_s1_readdata_from_sa => uart1_s1_readdata_from_sa
    );


  --the_pipeline_bridge, which is an e_ptf_instance
  the_pipeline_bridge : pipeline_bridge
    port map(
      m1_address => pipeline_bridge_m1_address,
      m1_burstcount => pipeline_bridge_m1_burstcount,
      m1_byteenable => pipeline_bridge_m1_byteenable,
      m1_chipselect => pipeline_bridge_m1_chipselect,
      m1_debugaccess => pipeline_bridge_m1_debugaccess,
      m1_read => pipeline_bridge_m1_read,
      m1_write => pipeline_bridge_m1_write,
      m1_writedata => pipeline_bridge_m1_writedata,
      s1_endofpacket => pipeline_bridge_s1_endofpacket,
      s1_readdata => pipeline_bridge_s1_readdata,
      s1_readdatavalid => pipeline_bridge_s1_readdatavalid,
      s1_waitrequest => pipeline_bridge_s1_waitrequest,
      clk => internal_pll_c0_out,
      m1_endofpacket => pipeline_bridge_m1_endofpacket,
      m1_readdata => pipeline_bridge_m1_readdata,
      m1_readdatavalid => pipeline_bridge_m1_readdatavalid,
      m1_waitrequest => pipeline_bridge_m1_waitrequest,
      reset_n => pipeline_bridge_s1_reset_n,
      s1_address => pipeline_bridge_s1_address,
      s1_arbiterlock => pipeline_bridge_s1_arbiterlock,
      s1_arbiterlock2 => pipeline_bridge_s1_arbiterlock2,
      s1_burstcount => pipeline_bridge_s1_burstcount,
      s1_byteenable => pipeline_bridge_s1_byteenable,
      s1_chipselect => pipeline_bridge_s1_chipselect,
      s1_debugaccess => pipeline_bridge_s1_debugaccess,
      s1_nativeaddress => pipeline_bridge_s1_nativeaddress,
      s1_read => pipeline_bridge_s1_read,
      s1_write => pipeline_bridge_s1_write,
      s1_writedata => pipeline_bridge_s1_writedata
    );


  --the_pll_s1, which is an e_instance
  the_pll_s1 : pll_s1_arbitrator
    port map(
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_granted_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_qualified_request_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_data_valid_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read_data_valid_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_requests_pll_s1,
      d1_pll_s1_end_xfer => d1_pll_s1_end_xfer,
      pll_s1_address => pll_s1_address,
      pll_s1_chipselect => pll_s1_chipselect,
      pll_s1_read => pll_s1_read,
      pll_s1_readdata_from_sa => pll_s1_readdata_from_sa,
      pll_s1_reset_n => pll_s1_reset_n,
      pll_s1_resetrequest_from_sa => pll_s1_resetrequest_from_sa,
      pll_s1_write => pll_s1_write,
      pll_s1_writedata => pll_s1_writedata,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_address_to_slave,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_nativeaddress => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_nativeaddress,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_read,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_write,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_writedata,
      clk => clk,
      pll_s1_readdata => pll_s1_readdata,
      pll_s1_resetrequest => pll_s1_resetrequest,
      reset_n => clk_reset_n
    );


  --pll_c0_out out_clk assignment, which is an e_assign
  internal_pll_c0_out <= out_clk_pll_c0;
  --pll_c1_out out_clk assignment, which is an e_assign
  pll_c1_out <= out_clk_pll_c1;
  --pll_c2_out out_clk assignment, which is an e_assign
  pll_c2_out <= out_clk_pll_c2;
  --the_pll, which is an e_ptf_instance
  the_pll : pll
    port map(
      c0 => out_clk_pll_c0,
      c1 => out_clk_pll_c1,
      c2 => out_clk_pll_c2,
      readdata => pll_s1_readdata,
      resetrequest => pll_s1_resetrequest,
      address => pll_s1_address,
      chipselect => pll_s1_chipselect,
      clk => clk,
      read => pll_s1_read,
      reset_n => pll_s1_reset_n,
      write => pll_s1_write,
      writedata => pll_s1_writedata
    );


  --the_reconfig_request_pio_s1, which is an e_instance
  the_reconfig_request_pio_s1 : reconfig_request_pio_s1_arbitrator
    port map(
      d1_reconfig_request_pio_s1_end_xfer => d1_reconfig_request_pio_s1_end_xfer,
      pipeline_bridge_m1_granted_reconfig_request_pio_s1 => pipeline_bridge_m1_granted_reconfig_request_pio_s1,
      pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1 => pipeline_bridge_m1_qualified_request_reconfig_request_pio_s1,
      pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1 => pipeline_bridge_m1_read_data_valid_reconfig_request_pio_s1,
      pipeline_bridge_m1_requests_reconfig_request_pio_s1 => pipeline_bridge_m1_requests_reconfig_request_pio_s1,
      reconfig_request_pio_s1_address => reconfig_request_pio_s1_address,
      reconfig_request_pio_s1_chipselect => reconfig_request_pio_s1_chipselect,
      reconfig_request_pio_s1_readdata_from_sa => reconfig_request_pio_s1_readdata_from_sa,
      reconfig_request_pio_s1_reset_n => reconfig_request_pio_s1_reset_n,
      reconfig_request_pio_s1_write_n => reconfig_request_pio_s1_write_n,
      reconfig_request_pio_s1_writedata => reconfig_request_pio_s1_writedata,
      clk => internal_pll_c0_out,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reconfig_request_pio_s1_readdata => reconfig_request_pio_s1_readdata,
      reset_n => pll_c0_out_reset_n
    );


  --the_reconfig_request_pio, which is an e_ptf_instance
  the_reconfig_request_pio : reconfig_request_pio
    port map(
      bidir_port => bidir_port_to_and_from_the_reconfig_request_pio,
      readdata => reconfig_request_pio_s1_readdata,
      address => reconfig_request_pio_s1_address,
      chipselect => reconfig_request_pio_s1_chipselect,
      clk => internal_pll_c0_out,
      reset_n => reconfig_request_pio_s1_reset_n,
      write_n => reconfig_request_pio_s1_write_n,
      writedata => reconfig_request_pio_s1_writedata
    );


  --the_seven_seg_pio_s1, which is an e_instance
  the_seven_seg_pio_s1 : seven_seg_pio_s1_arbitrator
    port map(
      d1_seven_seg_pio_s1_end_xfer => d1_seven_seg_pio_s1_end_xfer,
      pipeline_bridge_m1_granted_seven_seg_pio_s1 => pipeline_bridge_m1_granted_seven_seg_pio_s1,
      pipeline_bridge_m1_qualified_request_seven_seg_pio_s1 => pipeline_bridge_m1_qualified_request_seven_seg_pio_s1,
      pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1 => pipeline_bridge_m1_read_data_valid_seven_seg_pio_s1,
      pipeline_bridge_m1_requests_seven_seg_pio_s1 => pipeline_bridge_m1_requests_seven_seg_pio_s1,
      seven_seg_pio_s1_address => seven_seg_pio_s1_address,
      seven_seg_pio_s1_chipselect => seven_seg_pio_s1_chipselect,
      seven_seg_pio_s1_readdata_from_sa => seven_seg_pio_s1_readdata_from_sa,
      seven_seg_pio_s1_reset_n => seven_seg_pio_s1_reset_n,
      seven_seg_pio_s1_write_n => seven_seg_pio_s1_write_n,
      seven_seg_pio_s1_writedata => seven_seg_pio_s1_writedata,
      clk => internal_pll_c0_out,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n,
      seven_seg_pio_s1_readdata => seven_seg_pio_s1_readdata
    );


  --the_seven_seg_pio, which is an e_ptf_instance
  the_seven_seg_pio : seven_seg_pio
    port map(
      out_port => internal_out_port_from_the_seven_seg_pio,
      readdata => seven_seg_pio_s1_readdata,
      address => seven_seg_pio_s1_address,
      chipselect => seven_seg_pio_s1_chipselect,
      clk => internal_pll_c0_out,
      reset_n => seven_seg_pio_s1_reset_n,
      write_n => seven_seg_pio_s1_write_n,
      writedata => seven_seg_pio_s1_writedata
    );


  --the_sgdma_rx_csr, which is an e_instance
  the_sgdma_rx_csr : sgdma_rx_csr_arbitrator
    port map(
      d1_sgdma_rx_csr_end_xfer => d1_sgdma_rx_csr_end_xfer,
      pipeline_bridge_m1_granted_sgdma_rx_csr => pipeline_bridge_m1_granted_sgdma_rx_csr,
      pipeline_bridge_m1_qualified_request_sgdma_rx_csr => pipeline_bridge_m1_qualified_request_sgdma_rx_csr,
      pipeline_bridge_m1_read_data_valid_sgdma_rx_csr => pipeline_bridge_m1_read_data_valid_sgdma_rx_csr,
      pipeline_bridge_m1_requests_sgdma_rx_csr => pipeline_bridge_m1_requests_sgdma_rx_csr,
      sgdma_rx_csr_address => sgdma_rx_csr_address,
      sgdma_rx_csr_chipselect => sgdma_rx_csr_chipselect,
      sgdma_rx_csr_irq_from_sa => sgdma_rx_csr_irq_from_sa,
      sgdma_rx_csr_read => sgdma_rx_csr_read,
      sgdma_rx_csr_readdata_from_sa => sgdma_rx_csr_readdata_from_sa,
      sgdma_rx_csr_reset_n => sgdma_rx_csr_reset_n,
      sgdma_rx_csr_write => sgdma_rx_csr_write,
      sgdma_rx_csr_writedata => sgdma_rx_csr_writedata,
      clk => internal_pll_c0_out,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_csr_irq => sgdma_rx_csr_irq,
      sgdma_rx_csr_readdata => sgdma_rx_csr_readdata
    );


  --the_sgdma_rx_in, which is an e_instance
  the_sgdma_rx_in : sgdma_rx_in_arbitrator
    port map(
      sgdma_rx_in_data => sgdma_rx_in_data,
      sgdma_rx_in_empty => sgdma_rx_in_empty,
      sgdma_rx_in_endofpacket => sgdma_rx_in_endofpacket,
      sgdma_rx_in_error => sgdma_rx_in_error,
      sgdma_rx_in_ready_from_sa => sgdma_rx_in_ready_from_sa,
      sgdma_rx_in_startofpacket => sgdma_rx_in_startofpacket,
      sgdma_rx_in_valid => sgdma_rx_in_valid,
      clk => internal_pll_c0_out,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_in_ready => sgdma_rx_in_ready,
      tse_mac_receive_data => tse_mac_receive_data,
      tse_mac_receive_empty => tse_mac_receive_empty,
      tse_mac_receive_endofpacket => tse_mac_receive_endofpacket,
      tse_mac_receive_error => tse_mac_receive_error,
      tse_mac_receive_startofpacket => tse_mac_receive_startofpacket,
      tse_mac_receive_valid => tse_mac_receive_valid
    );


  --the_sgdma_rx_descriptor_read, which is an e_instance
  the_sgdma_rx_descriptor_read : sgdma_rx_descriptor_read_arbitrator
    port map(
      sgdma_rx_descriptor_read_address_to_slave => sgdma_rx_descriptor_read_address_to_slave,
      sgdma_rx_descriptor_read_latency_counter => sgdma_rx_descriptor_read_latency_counter,
      sgdma_rx_descriptor_read_readdata => sgdma_rx_descriptor_read_readdata,
      sgdma_rx_descriptor_read_readdatavalid => sgdma_rx_descriptor_read_readdatavalid,
      sgdma_rx_descriptor_read_waitrequest => sgdma_rx_descriptor_read_waitrequest,
      clk => internal_pll_c0_out,
      d1_descriptor_memory_s1_end_xfer => d1_descriptor_memory_s1_end_xfer,
      descriptor_memory_s1_readdata_from_sa => descriptor_memory_s1_readdata_from_sa,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_descriptor_read_address => sgdma_rx_descriptor_read_address,
      sgdma_rx_descriptor_read_granted_descriptor_memory_s1 => sgdma_rx_descriptor_read_granted_descriptor_memory_s1,
      sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1 => sgdma_rx_descriptor_read_qualified_request_descriptor_memory_s1,
      sgdma_rx_descriptor_read_read => sgdma_rx_descriptor_read_read,
      sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1 => sgdma_rx_descriptor_read_read_data_valid_descriptor_memory_s1,
      sgdma_rx_descriptor_read_requests_descriptor_memory_s1 => sgdma_rx_descriptor_read_requests_descriptor_memory_s1
    );


  --the_sgdma_rx_descriptor_write, which is an e_instance
  the_sgdma_rx_descriptor_write : sgdma_rx_descriptor_write_arbitrator
    port map(
      sgdma_rx_descriptor_write_address_to_slave => sgdma_rx_descriptor_write_address_to_slave,
      sgdma_rx_descriptor_write_waitrequest => sgdma_rx_descriptor_write_waitrequest,
      clk => internal_pll_c0_out,
      d1_descriptor_memory_s1_end_xfer => d1_descriptor_memory_s1_end_xfer,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_descriptor_write_address => sgdma_rx_descriptor_write_address,
      sgdma_rx_descriptor_write_granted_descriptor_memory_s1 => sgdma_rx_descriptor_write_granted_descriptor_memory_s1,
      sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1 => sgdma_rx_descriptor_write_qualified_request_descriptor_memory_s1,
      sgdma_rx_descriptor_write_requests_descriptor_memory_s1 => sgdma_rx_descriptor_write_requests_descriptor_memory_s1,
      sgdma_rx_descriptor_write_write => sgdma_rx_descriptor_write_write,
      sgdma_rx_descriptor_write_writedata => sgdma_rx_descriptor_write_writedata
    );


  --the_sgdma_rx_m_write, which is an e_instance
  the_sgdma_rx_m_write : sgdma_rx_m_write_arbitrator
    port map(
      sgdma_rx_m_write_address_to_slave => sgdma_rx_m_write_address_to_slave,
      sgdma_rx_m_write_waitrequest => sgdma_rx_m_write_waitrequest,
      clk => internal_pll_c0_out,
      d1_ddr_sdram_0_s1_end_xfer => d1_ddr_sdram_0_s1_end_xfer,
      d1_ext_ssram_bus_avalon_slave_end_xfer => d1_ext_ssram_bus_avalon_slave_end_xfer,
      d1_packet_memory_s2_end_xfer => d1_packet_memory_s2_end_xfer,
      ddr_sdram_0_s1_waitrequest_n_from_sa => ddr_sdram_0_s1_waitrequest_n_from_sa,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_m_write_address => sgdma_rx_m_write_address,
      sgdma_rx_m_write_byteenable => sgdma_rx_m_write_byteenable,
      sgdma_rx_m_write_granted_ddr_sdram_0_s1 => sgdma_rx_m_write_granted_ddr_sdram_0_s1,
      sgdma_rx_m_write_granted_ext_ssram_s1 => sgdma_rx_m_write_granted_ext_ssram_s1,
      sgdma_rx_m_write_granted_packet_memory_s2 => sgdma_rx_m_write_granted_packet_memory_s2,
      sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1 => sgdma_rx_m_write_qualified_request_ddr_sdram_0_s1,
      sgdma_rx_m_write_qualified_request_ext_ssram_s1 => sgdma_rx_m_write_qualified_request_ext_ssram_s1,
      sgdma_rx_m_write_qualified_request_packet_memory_s2 => sgdma_rx_m_write_qualified_request_packet_memory_s2,
      sgdma_rx_m_write_requests_ddr_sdram_0_s1 => sgdma_rx_m_write_requests_ddr_sdram_0_s1,
      sgdma_rx_m_write_requests_ext_ssram_s1 => sgdma_rx_m_write_requests_ext_ssram_s1,
      sgdma_rx_m_write_requests_packet_memory_s2 => sgdma_rx_m_write_requests_packet_memory_s2,
      sgdma_rx_m_write_write => sgdma_rx_m_write_write,
      sgdma_rx_m_write_writedata => sgdma_rx_m_write_writedata
    );


  --the_sgdma_rx, which is an e_ptf_instance
  the_sgdma_rx : sgdma_rx
    port map(
      csr_irq => sgdma_rx_csr_irq,
      csr_readdata => sgdma_rx_csr_readdata,
      descriptor_read_address => sgdma_rx_descriptor_read_address,
      descriptor_read_read => sgdma_rx_descriptor_read_read,
      descriptor_write_address => sgdma_rx_descriptor_write_address,
      descriptor_write_write => sgdma_rx_descriptor_write_write,
      descriptor_write_writedata => sgdma_rx_descriptor_write_writedata,
      in_ready => sgdma_rx_in_ready,
      m_write_address => sgdma_rx_m_write_address,
      m_write_byteenable => sgdma_rx_m_write_byteenable,
      m_write_write => sgdma_rx_m_write_write,
      m_write_writedata => sgdma_rx_m_write_writedata,
      clk => internal_pll_c0_out,
      csr_address => sgdma_rx_csr_address,
      csr_chipselect => sgdma_rx_csr_chipselect,
      csr_read => sgdma_rx_csr_read,
      csr_write => sgdma_rx_csr_write,
      csr_writedata => sgdma_rx_csr_writedata,
      descriptor_read_readdata => sgdma_rx_descriptor_read_readdata,
      descriptor_read_readdatavalid => sgdma_rx_descriptor_read_readdatavalid,
      descriptor_read_waitrequest => sgdma_rx_descriptor_read_waitrequest,
      descriptor_write_waitrequest => sgdma_rx_descriptor_write_waitrequest,
      in_data => sgdma_rx_in_data,
      in_empty => sgdma_rx_in_empty,
      in_endofpacket => sgdma_rx_in_endofpacket,
      in_error => sgdma_rx_in_error,
      in_startofpacket => sgdma_rx_in_startofpacket,
      in_valid => sgdma_rx_in_valid,
      m_write_waitrequest => sgdma_rx_m_write_waitrequest,
      system_reset_n => sgdma_rx_csr_reset_n
    );


  --the_sgdma_tx_csr, which is an e_instance
  the_sgdma_tx_csr : sgdma_tx_csr_arbitrator
    port map(
      d1_sgdma_tx_csr_end_xfer => d1_sgdma_tx_csr_end_xfer,
      pipeline_bridge_m1_granted_sgdma_tx_csr => pipeline_bridge_m1_granted_sgdma_tx_csr,
      pipeline_bridge_m1_qualified_request_sgdma_tx_csr => pipeline_bridge_m1_qualified_request_sgdma_tx_csr,
      pipeline_bridge_m1_read_data_valid_sgdma_tx_csr => pipeline_bridge_m1_read_data_valid_sgdma_tx_csr,
      pipeline_bridge_m1_requests_sgdma_tx_csr => pipeline_bridge_m1_requests_sgdma_tx_csr,
      sgdma_tx_csr_address => sgdma_tx_csr_address,
      sgdma_tx_csr_chipselect => sgdma_tx_csr_chipselect,
      sgdma_tx_csr_irq_from_sa => sgdma_tx_csr_irq_from_sa,
      sgdma_tx_csr_read => sgdma_tx_csr_read,
      sgdma_tx_csr_readdata_from_sa => sgdma_tx_csr_readdata_from_sa,
      sgdma_tx_csr_reset_n => sgdma_tx_csr_reset_n,
      sgdma_tx_csr_write => sgdma_tx_csr_write,
      sgdma_tx_csr_writedata => sgdma_tx_csr_writedata,
      clk => internal_pll_c0_out,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n,
      sgdma_tx_csr_irq => sgdma_tx_csr_irq,
      sgdma_tx_csr_readdata => sgdma_tx_csr_readdata
    );


  --the_sgdma_tx_descriptor_read, which is an e_instance
  the_sgdma_tx_descriptor_read : sgdma_tx_descriptor_read_arbitrator
    port map(
      sgdma_tx_descriptor_read_address_to_slave => sgdma_tx_descriptor_read_address_to_slave,
      sgdma_tx_descriptor_read_latency_counter => sgdma_tx_descriptor_read_latency_counter,
      sgdma_tx_descriptor_read_readdata => sgdma_tx_descriptor_read_readdata,
      sgdma_tx_descriptor_read_readdatavalid => sgdma_tx_descriptor_read_readdatavalid,
      sgdma_tx_descriptor_read_waitrequest => sgdma_tx_descriptor_read_waitrequest,
      clk => internal_pll_c0_out,
      d1_descriptor_memory_s1_end_xfer => d1_descriptor_memory_s1_end_xfer,
      descriptor_memory_s1_readdata_from_sa => descriptor_memory_s1_readdata_from_sa,
      reset_n => pll_c0_out_reset_n,
      sgdma_tx_descriptor_read_address => sgdma_tx_descriptor_read_address,
      sgdma_tx_descriptor_read_granted_descriptor_memory_s1 => sgdma_tx_descriptor_read_granted_descriptor_memory_s1,
      sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1 => sgdma_tx_descriptor_read_qualified_request_descriptor_memory_s1,
      sgdma_tx_descriptor_read_read => sgdma_tx_descriptor_read_read,
      sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1 => sgdma_tx_descriptor_read_read_data_valid_descriptor_memory_s1,
      sgdma_tx_descriptor_read_requests_descriptor_memory_s1 => sgdma_tx_descriptor_read_requests_descriptor_memory_s1
    );


  --the_sgdma_tx_descriptor_write, which is an e_instance
  the_sgdma_tx_descriptor_write : sgdma_tx_descriptor_write_arbitrator
    port map(
      sgdma_tx_descriptor_write_address_to_slave => sgdma_tx_descriptor_write_address_to_slave,
      sgdma_tx_descriptor_write_waitrequest => sgdma_tx_descriptor_write_waitrequest,
      clk => internal_pll_c0_out,
      d1_descriptor_memory_s1_end_xfer => d1_descriptor_memory_s1_end_xfer,
      reset_n => pll_c0_out_reset_n,
      sgdma_tx_descriptor_write_address => sgdma_tx_descriptor_write_address,
      sgdma_tx_descriptor_write_granted_descriptor_memory_s1 => sgdma_tx_descriptor_write_granted_descriptor_memory_s1,
      sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1 => sgdma_tx_descriptor_write_qualified_request_descriptor_memory_s1,
      sgdma_tx_descriptor_write_requests_descriptor_memory_s1 => sgdma_tx_descriptor_write_requests_descriptor_memory_s1,
      sgdma_tx_descriptor_write_write => sgdma_tx_descriptor_write_write,
      sgdma_tx_descriptor_write_writedata => sgdma_tx_descriptor_write_writedata
    );


  --the_sgdma_tx_m_read, which is an e_instance
  the_sgdma_tx_m_read : sgdma_tx_m_read_arbitrator
    port map(
      sgdma_tx_m_read_address_to_slave => sgdma_tx_m_read_address_to_slave,
      sgdma_tx_m_read_latency_counter => sgdma_tx_m_read_latency_counter,
      sgdma_tx_m_read_readdata => sgdma_tx_m_read_readdata,
      sgdma_tx_m_read_readdatavalid => sgdma_tx_m_read_readdatavalid,
      sgdma_tx_m_read_waitrequest => sgdma_tx_m_read_waitrequest,
      clk => internal_pll_c0_out,
      d1_ddr_sdram_0_s1_end_xfer => d1_ddr_sdram_0_s1_end_xfer,
      d1_ext_ssram_bus_avalon_slave_end_xfer => d1_ext_ssram_bus_avalon_slave_end_xfer,
      d1_packet_memory_s2_end_xfer => d1_packet_memory_s2_end_xfer,
      ddr_sdram_0_s1_readdata_from_sa => ddr_sdram_0_s1_readdata_from_sa,
      ddr_sdram_0_s1_waitrequest_n_from_sa => ddr_sdram_0_s1_waitrequest_n_from_sa,
      incoming_ext_ssram_bus_data => incoming_ext_ssram_bus_data,
      packet_memory_s2_readdata_from_sa => packet_memory_s2_readdata_from_sa,
      reset_n => pll_c0_out_reset_n,
      sgdma_tx_m_read_address => sgdma_tx_m_read_address,
      sgdma_tx_m_read_granted_ddr_sdram_0_s1 => sgdma_tx_m_read_granted_ddr_sdram_0_s1,
      sgdma_tx_m_read_granted_ext_ssram_s1 => sgdma_tx_m_read_granted_ext_ssram_s1,
      sgdma_tx_m_read_granted_packet_memory_s2 => sgdma_tx_m_read_granted_packet_memory_s2,
      sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1 => sgdma_tx_m_read_qualified_request_ddr_sdram_0_s1,
      sgdma_tx_m_read_qualified_request_ext_ssram_s1 => sgdma_tx_m_read_qualified_request_ext_ssram_s1,
      sgdma_tx_m_read_qualified_request_packet_memory_s2 => sgdma_tx_m_read_qualified_request_packet_memory_s2,
      sgdma_tx_m_read_read => sgdma_tx_m_read_read,
      sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1 => sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1,
      sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register => sgdma_tx_m_read_read_data_valid_ddr_sdram_0_s1_shift_register,
      sgdma_tx_m_read_read_data_valid_ext_ssram_s1 => sgdma_tx_m_read_read_data_valid_ext_ssram_s1,
      sgdma_tx_m_read_read_data_valid_packet_memory_s2 => sgdma_tx_m_read_read_data_valid_packet_memory_s2,
      sgdma_tx_m_read_requests_ddr_sdram_0_s1 => sgdma_tx_m_read_requests_ddr_sdram_0_s1,
      sgdma_tx_m_read_requests_ext_ssram_s1 => sgdma_tx_m_read_requests_ext_ssram_s1,
      sgdma_tx_m_read_requests_packet_memory_s2 => sgdma_tx_m_read_requests_packet_memory_s2
    );


  --the_sgdma_tx_out, which is an e_instance
  the_sgdma_tx_out : sgdma_tx_out_arbitrator
    port map(
      sgdma_tx_out_ready => sgdma_tx_out_ready,
      clk => internal_pll_c0_out,
      reset_n => pll_c0_out_reset_n,
      sgdma_tx_out_data => sgdma_tx_out_data,
      sgdma_tx_out_empty => sgdma_tx_out_empty,
      sgdma_tx_out_endofpacket => sgdma_tx_out_endofpacket,
      sgdma_tx_out_error => sgdma_tx_out_error,
      sgdma_tx_out_startofpacket => sgdma_tx_out_startofpacket,
      sgdma_tx_out_valid => sgdma_tx_out_valid,
      tse_mac_transmit_ready_from_sa => tse_mac_transmit_ready_from_sa
    );


  --the_sgdma_tx, which is an e_ptf_instance
  the_sgdma_tx : sgdma_tx
    port map(
      csr_irq => sgdma_tx_csr_irq,
      csr_readdata => sgdma_tx_csr_readdata,
      descriptor_read_address => sgdma_tx_descriptor_read_address,
      descriptor_read_read => sgdma_tx_descriptor_read_read,
      descriptor_write_address => sgdma_tx_descriptor_write_address,
      descriptor_write_write => sgdma_tx_descriptor_write_write,
      descriptor_write_writedata => sgdma_tx_descriptor_write_writedata,
      m_read_address => sgdma_tx_m_read_address,
      m_read_read => sgdma_tx_m_read_read,
      out_data => sgdma_tx_out_data,
      out_empty => sgdma_tx_out_empty,
      out_endofpacket => sgdma_tx_out_endofpacket,
      out_error => sgdma_tx_out_error,
      out_startofpacket => sgdma_tx_out_startofpacket,
      out_valid => sgdma_tx_out_valid,
      clk => internal_pll_c0_out,
      csr_address => sgdma_tx_csr_address,
      csr_chipselect => sgdma_tx_csr_chipselect,
      csr_read => sgdma_tx_csr_read,
      csr_write => sgdma_tx_csr_write,
      csr_writedata => sgdma_tx_csr_writedata,
      descriptor_read_readdata => sgdma_tx_descriptor_read_readdata,
      descriptor_read_readdatavalid => sgdma_tx_descriptor_read_readdatavalid,
      descriptor_read_waitrequest => sgdma_tx_descriptor_read_waitrequest,
      descriptor_write_waitrequest => sgdma_tx_descriptor_write_waitrequest,
      m_read_readdata => sgdma_tx_m_read_readdata,
      m_read_readdatavalid => sgdma_tx_m_read_readdatavalid,
      m_read_waitrequest => sgdma_tx_m_read_waitrequest,
      out_ready => sgdma_tx_out_ready,
      system_reset_n => sgdma_tx_csr_reset_n
    );


  --the_sys_clk_timer_s1, which is an e_instance
  the_sys_clk_timer_s1 : sys_clk_timer_s1_arbitrator
    port map(
      d1_sys_clk_timer_s1_end_xfer => d1_sys_clk_timer_s1_end_xfer,
      pipeline_bridge_m1_granted_sys_clk_timer_s1 => pipeline_bridge_m1_granted_sys_clk_timer_s1,
      pipeline_bridge_m1_qualified_request_sys_clk_timer_s1 => pipeline_bridge_m1_qualified_request_sys_clk_timer_s1,
      pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1 => pipeline_bridge_m1_read_data_valid_sys_clk_timer_s1,
      pipeline_bridge_m1_requests_sys_clk_timer_s1 => pipeline_bridge_m1_requests_sys_clk_timer_s1,
      sys_clk_timer_s1_address => sys_clk_timer_s1_address,
      sys_clk_timer_s1_chipselect => sys_clk_timer_s1_chipselect,
      sys_clk_timer_s1_irq_from_sa => sys_clk_timer_s1_irq_from_sa,
      sys_clk_timer_s1_readdata_from_sa => sys_clk_timer_s1_readdata_from_sa,
      sys_clk_timer_s1_reset_n => sys_clk_timer_s1_reset_n,
      sys_clk_timer_s1_write_n => sys_clk_timer_s1_write_n,
      sys_clk_timer_s1_writedata => sys_clk_timer_s1_writedata,
      clk => internal_pll_c0_out,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n,
      sys_clk_timer_s1_irq => sys_clk_timer_s1_irq,
      sys_clk_timer_s1_readdata => sys_clk_timer_s1_readdata
    );


  --the_sys_clk_timer, which is an e_ptf_instance
  the_sys_clk_timer : sys_clk_timer
    port map(
      irq => sys_clk_timer_s1_irq,
      readdata => sys_clk_timer_s1_readdata,
      address => sys_clk_timer_s1_address,
      chipselect => sys_clk_timer_s1_chipselect,
      clk => internal_pll_c0_out,
      reset_n => sys_clk_timer_s1_reset_n,
      write_n => sys_clk_timer_s1_write_n,
      writedata => sys_clk_timer_s1_writedata
    );


  --the_tse_mac_control_port, which is an e_instance
  the_tse_mac_control_port : tse_mac_control_port_arbitrator
    port map(
      cpu_data_master_granted_tse_mac_control_port => cpu_data_master_granted_tse_mac_control_port,
      cpu_data_master_qualified_request_tse_mac_control_port => cpu_data_master_qualified_request_tse_mac_control_port,
      cpu_data_master_read_data_valid_tse_mac_control_port => cpu_data_master_read_data_valid_tse_mac_control_port,
      cpu_data_master_requests_tse_mac_control_port => cpu_data_master_requests_tse_mac_control_port,
      d1_tse_mac_control_port_end_xfer => d1_tse_mac_control_port_end_xfer,
      tse_mac_control_port_address => tse_mac_control_port_address,
      tse_mac_control_port_read => tse_mac_control_port_read,
      tse_mac_control_port_readdata_from_sa => tse_mac_control_port_readdata_from_sa,
      tse_mac_control_port_reset => tse_mac_control_port_reset,
      tse_mac_control_port_waitrequest_from_sa => tse_mac_control_port_waitrequest_from_sa,
      tse_mac_control_port_write => tse_mac_control_port_write,
      tse_mac_control_port_writedata => tse_mac_control_port_writedata,
      clk => internal_pll_c0_out,
      cpu_data_master_address_to_slave => cpu_data_master_address_to_slave,
      cpu_data_master_latency_counter => cpu_data_master_latency_counter,
      cpu_data_master_read => cpu_data_master_read,
      cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register => cpu_data_master_read_data_valid_ddr_sdram_0_s1_shift_register,
      cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register => cpu_data_master_read_data_valid_pipeline_bridge_s1_shift_register,
      cpu_data_master_write => cpu_data_master_write,
      cpu_data_master_writedata => cpu_data_master_writedata,
      reset_n => pll_c0_out_reset_n,
      tse_mac_control_port_readdata => tse_mac_control_port_readdata,
      tse_mac_control_port_waitrequest => tse_mac_control_port_waitrequest
    );


  --the_tse_mac_transmit, which is an e_instance
  the_tse_mac_transmit : tse_mac_transmit_arbitrator
    port map(
      tse_mac_transmit_data => tse_mac_transmit_data,
      tse_mac_transmit_empty => tse_mac_transmit_empty,
      tse_mac_transmit_endofpacket => tse_mac_transmit_endofpacket,
      tse_mac_transmit_error => tse_mac_transmit_error,
      tse_mac_transmit_ready_from_sa => tse_mac_transmit_ready_from_sa,
      tse_mac_transmit_startofpacket => tse_mac_transmit_startofpacket,
      tse_mac_transmit_valid => tse_mac_transmit_valid,
      clk => internal_pll_c0_out,
      reset_n => pll_c0_out_reset_n,
      sgdma_tx_out_data => sgdma_tx_out_data,
      sgdma_tx_out_empty => sgdma_tx_out_empty,
      sgdma_tx_out_endofpacket => sgdma_tx_out_endofpacket,
      sgdma_tx_out_error => sgdma_tx_out_error,
      sgdma_tx_out_startofpacket => sgdma_tx_out_startofpacket,
      sgdma_tx_out_valid => sgdma_tx_out_valid,
      tse_mac_transmit_ready => tse_mac_transmit_ready
    );


  --the_tse_mac_receive, which is an e_instance
  the_tse_mac_receive : tse_mac_receive_arbitrator
    port map(
      tse_mac_receive_ready => tse_mac_receive_ready,
      clk => internal_pll_c0_out,
      reset_n => pll_c0_out_reset_n,
      sgdma_rx_in_ready_from_sa => sgdma_rx_in_ready_from_sa,
      tse_mac_receive_data => tse_mac_receive_data,
      tse_mac_receive_empty => tse_mac_receive_empty,
      tse_mac_receive_endofpacket => tse_mac_receive_endofpacket,
      tse_mac_receive_error => tse_mac_receive_error,
      tse_mac_receive_startofpacket => tse_mac_receive_startofpacket,
      tse_mac_receive_valid => tse_mac_receive_valid
    );


  --the_tse_mac, which is an e_ptf_instance
  the_tse_mac : tse_mac
    port map(
      ena_10 => internal_ena_10_from_the_tse_mac,
      eth_mode => internal_eth_mode_from_the_tse_mac,
      ff_rx_data => tse_mac_receive_data,
      ff_rx_dval => tse_mac_receive_valid,
      ff_rx_eop => tse_mac_receive_endofpacket,
      ff_rx_mod => tse_mac_receive_empty,
      ff_rx_sop => tse_mac_receive_startofpacket,
      ff_tx_rdy => tse_mac_transmit_ready,
      gm_tx_d => internal_gm_tx_d_from_the_tse_mac,
      gm_tx_en => internal_gm_tx_en_from_the_tse_mac,
      gm_tx_err => internal_gm_tx_err_from_the_tse_mac,
      m_tx_d => internal_m_tx_d_from_the_tse_mac,
      m_tx_en => internal_m_tx_en_from_the_tse_mac,
      m_tx_err => internal_m_tx_err_from_the_tse_mac,
      mdc => internal_mdc_from_the_tse_mac,
      mdio_oen => internal_mdio_oen_from_the_tse_mac,
      mdio_out => internal_mdio_out_from_the_tse_mac,
      readdata => tse_mac_control_port_readdata,
      rx_err => tse_mac_receive_error,
      waitrequest => tse_mac_control_port_waitrequest,
      address => tse_mac_control_port_address,
      clk => internal_pll_c0_out,
      ff_rx_clk => internal_pll_c0_out,
      ff_rx_rdy => tse_mac_receive_ready,
      ff_tx_clk => internal_pll_c0_out,
      ff_tx_data => tse_mac_transmit_data,
      ff_tx_eop => tse_mac_transmit_endofpacket,
      ff_tx_err => tse_mac_transmit_error,
      ff_tx_mod => tse_mac_transmit_empty,
      ff_tx_sop => tse_mac_transmit_startofpacket,
      ff_tx_wren => tse_mac_transmit_valid,
      gm_rx_d => gm_rx_d_to_the_tse_mac,
      gm_rx_dv => gm_rx_dv_to_the_tse_mac,
      gm_rx_err => gm_rx_err_to_the_tse_mac,
      m_rx_col => m_rx_col_to_the_tse_mac,
      m_rx_crs => m_rx_crs_to_the_tse_mac,
      m_rx_d => m_rx_d_to_the_tse_mac,
      m_rx_en => m_rx_en_to_the_tse_mac,
      m_rx_err => m_rx_err_to_the_tse_mac,
      mdio_in => mdio_in_to_the_tse_mac,
      read => tse_mac_control_port_read,
      reset => tse_mac_control_port_reset,
      rx_clk => rx_clk_to_the_tse_mac,
      set_10 => set_10_to_the_tse_mac,
      set_1000 => set_1000_to_the_tse_mac,
      tx_clk => tx_clk_to_the_tse_mac,
      write => tse_mac_control_port_write,
      writedata => tse_mac_control_port_writedata
    );


  --the_tse_pll_s1, which is an e_instance
  the_tse_pll_s1 : tse_pll_s1_arbitrator
    port map(
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_granted_tse_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_qualified_request_tse_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_data_valid_tse_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read_data_valid_tse_pll_s1,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1 => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_requests_tse_pll_s1,
      d1_tse_pll_s1_end_xfer => d1_tse_pll_s1_end_xfer,
      tse_pll_s1_address => tse_pll_s1_address,
      tse_pll_s1_chipselect => tse_pll_s1_chipselect,
      tse_pll_s1_read => tse_pll_s1_read,
      tse_pll_s1_readdata_from_sa => tse_pll_s1_readdata_from_sa,
      tse_pll_s1_reset_n => tse_pll_s1_reset_n,
      tse_pll_s1_resetrequest_from_sa => tse_pll_s1_resetrequest_from_sa,
      tse_pll_s1_write => tse_pll_s1_write,
      tse_pll_s1_writedata => tse_pll_s1_writedata,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_address_to_slave,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_nativeaddress => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_nativeaddress,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_read,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_write,
      NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata => NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_writedata,
      clk => clk_to_tse_pll,
      reset_n => clk_to_tse_pll_reset_n,
      tse_pll_s1_readdata => tse_pll_s1_readdata,
      tse_pll_s1_resetrequest => tse_pll_s1_resetrequest
    );


  --tse_pll_c0_out out_clk assignment, which is an e_assign
  tse_pll_c0_out <= out_clk_tse_pll_c0;
  --the_tse_pll, which is an e_ptf_instance
  the_tse_pll : tse_pll
    port map(
      c0 => out_clk_tse_pll_c0,
      readdata => tse_pll_s1_readdata,
      resetrequest => tse_pll_s1_resetrequest,
      address => tse_pll_s1_address,
      chipselect => tse_pll_s1_chipselect,
      clk => clk_to_tse_pll,
      read => tse_pll_s1_read,
      reset_n => tse_pll_s1_reset_n,
      write => tse_pll_s1_write,
      writedata => tse_pll_s1_writedata
    );


  --the_uart1_s1, which is an e_instance
  the_uart1_s1 : uart1_s1_arbitrator
    port map(
      d1_uart1_s1_end_xfer => d1_uart1_s1_end_xfer,
      pipeline_bridge_m1_granted_uart1_s1 => pipeline_bridge_m1_granted_uart1_s1,
      pipeline_bridge_m1_qualified_request_uart1_s1 => pipeline_bridge_m1_qualified_request_uart1_s1,
      pipeline_bridge_m1_read_data_valid_uart1_s1 => pipeline_bridge_m1_read_data_valid_uart1_s1,
      pipeline_bridge_m1_requests_uart1_s1 => pipeline_bridge_m1_requests_uart1_s1,
      uart1_s1_address => uart1_s1_address,
      uart1_s1_begintransfer => uart1_s1_begintransfer,
      uart1_s1_chipselect => uart1_s1_chipselect,
      uart1_s1_dataavailable_from_sa => uart1_s1_dataavailable_from_sa,
      uart1_s1_irq_from_sa => uart1_s1_irq_from_sa,
      uart1_s1_read_n => uart1_s1_read_n,
      uart1_s1_readdata_from_sa => uart1_s1_readdata_from_sa,
      uart1_s1_readyfordata_from_sa => uart1_s1_readyfordata_from_sa,
      uart1_s1_reset_n => uart1_s1_reset_n,
      uart1_s1_write_n => uart1_s1_write_n,
      uart1_s1_writedata => uart1_s1_writedata,
      clk => internal_pll_c0_out,
      pipeline_bridge_m1_address_to_slave => pipeline_bridge_m1_address_to_slave,
      pipeline_bridge_m1_burstcount => pipeline_bridge_m1_burstcount,
      pipeline_bridge_m1_chipselect => pipeline_bridge_m1_chipselect,
      pipeline_bridge_m1_latency_counter => pipeline_bridge_m1_latency_counter,
      pipeline_bridge_m1_read => pipeline_bridge_m1_read,
      pipeline_bridge_m1_write => pipeline_bridge_m1_write,
      pipeline_bridge_m1_writedata => pipeline_bridge_m1_writedata,
      reset_n => pll_c0_out_reset_n,
      uart1_s1_dataavailable => uart1_s1_dataavailable,
      uart1_s1_irq => uart1_s1_irq,
      uart1_s1_readdata => uart1_s1_readdata,
      uart1_s1_readyfordata => uart1_s1_readyfordata
    );


  --the_uart1, which is an e_ptf_instance
  the_uart1 : uart1
    port map(
      dataavailable => uart1_s1_dataavailable,
      irq => uart1_s1_irq,
      readdata => uart1_s1_readdata,
      readyfordata => uart1_s1_readyfordata,
      txd => internal_txd_from_the_uart1,
      address => uart1_s1_address,
      begintransfer => uart1_s1_begintransfer,
      chipselect => uart1_s1_chipselect,
      clk => internal_pll_c0_out,
      read_n => uart1_s1_read_n,
      reset_n => uart1_s1_reset_n,
      rxd => rxd_to_the_uart1,
      write_n => uart1_s1_write_n,
      writedata => uart1_s1_writedata
    );


  --reset is asserted asynchronously and deasserted synchronously
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_pll_c0_out_domain_synch : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_pll_c0_out_domain_synch_module
    port map(
      data_out => pll_c0_out_reset_n,
      clk => internal_pll_c0_out,
      data_in => module_input15,
      reset_n => reset_n_sources
    );

  module_input15 <= std_logic'('1');

  --reset sources mux, which is an e_mux
  reset_n_sources <= Vector_To_Std_Logic(NOT (((((((((((std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(NOT reset_n))) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(cpu_jtag_debug_module_resetrequest_from_sa)))) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pll_s1_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(pll_s1_resetrequest_from_sa)))) OR std_logic_vector'("00000000000000000000000000000000")) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_pll_s1_resetrequest_from_sa)))) OR (std_logic_vector'("0000000000000000000000000000000") & (A_TOSTDLOGICVECTOR(tse_pll_s1_resetrequest_from_sa))))));
  --reset is asserted asynchronously and deasserted synchronously
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_domain_synch : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_domain_synch_module
    port map(
      data_out => clk_reset_n,
      clk => clk,
      data_in => module_input16,
      reset_n => reset_n_sources
    );

  module_input16 <= std_logic'('1');

  --reset is asserted asynchronously and deasserted synchronously
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_to_tse_pll_domain_synch : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_reset_clk_to_tse_pll_domain_synch_module
    port map(
      data_out => clk_to_tse_pll_reset_n,
      clk => clk_to_tse_pll,
      data_in => module_input17,
      reset_n => reset_n_sources
    );

  module_input17 <= std_logic'('1');

  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_endofpacket <= std_logic'('0');
  --NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_endofpacket of type endofpacket does not connect to anything so wire it to default (0)
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_endofpacket <= std_logic'('0');
  --vhdl renameroo for output signals
  LCD_E_from_the_lcd_display <= internal_LCD_E_from_the_lcd_display;
  --vhdl renameroo for output signals
  LCD_RS_from_the_lcd_display <= internal_LCD_RS_from_the_lcd_display;
  --vhdl renameroo for output signals
  LCD_RW_from_the_lcd_display <= internal_LCD_RW_from_the_lcd_display;
  --vhdl renameroo for output signals
  adsc_n_to_the_ext_ssram <= internal_adsc_n_to_the_ext_ssram;
  --vhdl renameroo for output signals
  bw_n_to_the_ext_ssram <= internal_bw_n_to_the_ext_ssram;
  --vhdl renameroo for output signals
  bwe_n_to_the_ext_ssram <= internal_bwe_n_to_the_ext_ssram;
  --vhdl renameroo for output signals
  chipenable1_n_to_the_ext_ssram <= internal_chipenable1_n_to_the_ext_ssram;
  --vhdl renameroo for output signals
  clk_to_sdram_from_the_ddr_sdram_0 <= internal_clk_to_sdram_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  clk_to_sdram_n_from_the_ddr_sdram_0 <= internal_clk_to_sdram_n_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  ddr_a_from_the_ddr_sdram_0 <= internal_ddr_a_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  ddr_ba_from_the_ddr_sdram_0 <= internal_ddr_ba_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  ddr_cas_n_from_the_ddr_sdram_0 <= internal_ddr_cas_n_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  ddr_cke_from_the_ddr_sdram_0 <= internal_ddr_cke_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  ddr_cs_n_from_the_ddr_sdram_0 <= internal_ddr_cs_n_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  ddr_dm_from_the_ddr_sdram_0 <= internal_ddr_dm_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  ddr_ras_n_from_the_ddr_sdram_0 <= internal_ddr_ras_n_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  ddr_we_n_from_the_ddr_sdram_0 <= internal_ddr_we_n_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  ena_10_from_the_tse_mac <= internal_ena_10_from_the_tse_mac;
  --vhdl renameroo for output signals
  eth_mode_from_the_tse_mac <= internal_eth_mode_from_the_tse_mac;
  --vhdl renameroo for output signals
  ext_flash_enet_bus_address <= internal_ext_flash_enet_bus_address;
  --vhdl renameroo for output signals
  ext_ssram_bus_address <= internal_ext_ssram_bus_address;
  --vhdl renameroo for output signals
  gm_tx_d_from_the_tse_mac <= internal_gm_tx_d_from_the_tse_mac;
  --vhdl renameroo for output signals
  gm_tx_en_from_the_tse_mac <= internal_gm_tx_en_from_the_tse_mac;
  --vhdl renameroo for output signals
  gm_tx_err_from_the_tse_mac <= internal_gm_tx_err_from_the_tse_mac;
  --vhdl renameroo for output signals
  jtag_debug_offchip_trace_clk_from_the_cpu <= internal_jtag_debug_offchip_trace_clk_from_the_cpu;
  --vhdl renameroo for output signals
  jtag_debug_offchip_trace_data_from_the_cpu <= internal_jtag_debug_offchip_trace_data_from_the_cpu;
  --vhdl renameroo for output signals
  jtag_debug_trigout_from_the_cpu <= internal_jtag_debug_trigout_from_the_cpu;
  --vhdl renameroo for output signals
  m_tx_d_from_the_tse_mac <= internal_m_tx_d_from_the_tse_mac;
  --vhdl renameroo for output signals
  m_tx_en_from_the_tse_mac <= internal_m_tx_en_from_the_tse_mac;
  --vhdl renameroo for output signals
  m_tx_err_from_the_tse_mac <= internal_m_tx_err_from_the_tse_mac;
  --vhdl renameroo for output signals
  mdc_from_the_tse_mac <= internal_mdc_from_the_tse_mac;
  --vhdl renameroo for output signals
  mdio_oen_from_the_tse_mac <= internal_mdio_oen_from_the_tse_mac;
  --vhdl renameroo for output signals
  mdio_out_from_the_tse_mac <= internal_mdio_out_from_the_tse_mac;
  --vhdl renameroo for output signals
  out_port_from_the_led_pio <= internal_out_port_from_the_led_pio;
  --vhdl renameroo for output signals
  out_port_from_the_seven_seg_pio <= internal_out_port_from_the_seven_seg_pio;
  --vhdl renameroo for output signals
  outputenable_n_to_the_ext_ssram <= internal_outputenable_n_to_the_ext_ssram;
  --vhdl renameroo for output signals
  pll_c0_out <= internal_pll_c0_out;
  --vhdl renameroo for output signals
  read_n_to_the_ext_flash <= internal_read_n_to_the_ext_flash;
  --vhdl renameroo for output signals
  select_n_to_the_ext_flash <= internal_select_n_to_the_ext_flash;
  --vhdl renameroo for output signals
  stratix_dll_control_from_the_ddr_sdram_0 <= internal_stratix_dll_control_from_the_ddr_sdram_0;
  --vhdl renameroo for output signals
  txd_from_the_uart1 <= internal_txd_from_the_uart1;
  --vhdl renameroo for output signals
  write_n_to_the_ext_flash <= internal_write_n_to_the_ext_flash;

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ext_flash_lane0_module is 
        port (
              -- inputs:
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ext_flash_lane0_module;


architecture europa of ext_flash_lane0_module is
              signal internal_q :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 16777215 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, rdaddress) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (23 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "ext_flash.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 16777216) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rdaddress)));
      


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity ext_flash_lane0_module is 
--        port (
--              
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity ext_flash_lane0_module;
--
--
--architecture europa of ext_flash_lane0_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal internal_q :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 16777215 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
--
--begin
--
--  process (rdaddress)
--  begin
--      read_address <= rdaddress;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "ext_flash.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "UNREGISTERED",
--      lpm_rdaddress_control => "UNREGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 24,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ext_flash is 
        port (
              -- inputs:
                 signal address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                 signal read_n : IN STD_LOGIC;
                 signal select_n : IN STD_LOGIC;
                 signal write_n : IN STD_LOGIC;

              -- outputs:
                 signal data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ext_flash;


architecture europa of ext_flash is
--synthesis translate_off
component ext_flash_lane0_module is 
           port (
                 -- inputs:
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ext_flash_lane0_module;

--synthesis translate_on
                signal data_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal logic_vector_gasket :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal module_input18 :  STD_LOGIC;
                signal module_input19 :  STD_LOGIC;
                signal q_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);

begin

  --s1, which is an e_ptf_slave
--synthesis translate_off
    logic_vector_gasket <= data;
    data_0 <= logic_vector_gasket(7 DOWNTO 0);
    --ext_flash_lane0, which is an e_ram
    ext_flash_lane0 : ext_flash_lane0_module
      port map(
        q => q_0,
        data => data_0,
        rdaddress => address,
        rdclken => module_input18,
        wraddress => address,
        wrclock => write_n,
        wren => module_input19
      );

    module_input18 <= std_logic'('1');
    module_input19 <= NOT select_n;

    data <= A_WE_StdLogicVector((std_logic'(((NOT select_n AND NOT read_n))) = '1'), q_0, A_REP(std_logic'('Z'), 8));
--synthesis translate_on

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ext_ssram_lane0_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ext_ssram_lane0_module;


architecture europa of ext_ssram_lane0_module is
              signal d1_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
              signal d2_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
              signal internal_q1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 524287 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, clk) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;
    VARIABLE rd_address_internal : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    VARIABLE d1_rdaddress : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    VARIABLE d2_rdaddress : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "ext_ssram_lane0.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 524288) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rd_address_internal)));
      
			 IF clk'event AND clk = '1' AND rdclken = '1' THEN
                            rd_address_internal := d2_rdaddress;
                            d2_rdaddress := d1_rdaddress;
                            d1_rdaddress := rdaddress;

                         END IF;
                        


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity ext_ssram_lane0_module is 
--        port (
--              
--                 signal clk : IN STD_LOGIC;
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal reset_n : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity ext_ssram_lane0_module;
--
--
--architecture europa of ext_ssram_lane0_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal rdclock : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal d1_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--                signal d2_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--                signal internal_q1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 524287 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--
--begin
--
--  process (clk, reset_n)
--  begin
--    if reset_n = '0' then
--      read_address <= std_logic_vector'("0000000000000000000");
--      read_address <= std_logic_vector'("0000000000000000000");
--    elsif clk'event and clk = '1' then
--      if std_logic'(rdclken) = '1' then 
--        read_address <= rdaddress;
--      end if;
--    end if;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "ext_ssram_lane0.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "REGISTERED",
--      lpm_rdaddress_control => "REGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 19,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q1,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            rdclock => clk,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q1;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ext_ssram_lane1_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ext_ssram_lane1_module;


architecture europa of ext_ssram_lane1_module is
              signal d1_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
              signal d2_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
              signal internal_q2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 524287 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, clk) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;
    VARIABLE rd_address_internal : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    VARIABLE d1_rdaddress : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    VARIABLE d2_rdaddress : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "ext_ssram_lane1.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 524288) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rd_address_internal)));
      
			 IF clk'event AND clk = '1' AND rdclken = '1' THEN
                            rd_address_internal := d2_rdaddress;
                            d2_rdaddress := d1_rdaddress;
                            d1_rdaddress := rdaddress;

                         END IF;
                        


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity ext_ssram_lane1_module is 
--        port (
--              
--                 signal clk : IN STD_LOGIC;
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal reset_n : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity ext_ssram_lane1_module;
--
--
--architecture europa of ext_ssram_lane1_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal rdclock : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal d1_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--                signal d2_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--                signal internal_q2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 524287 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--
--begin
--
--  process (clk, reset_n)
--  begin
--    if reset_n = '0' then
--      read_address <= std_logic_vector'("0000000000000000000");
--      read_address <= std_logic_vector'("0000000000000000000");
--    elsif clk'event and clk = '1' then
--      if std_logic'(rdclken) = '1' then 
--        read_address <= rdaddress;
--      end if;
--    end if;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "ext_ssram_lane1.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "REGISTERED",
--      lpm_rdaddress_control => "REGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 19,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q2,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            rdclock => clk,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q2;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ext_ssram_lane2_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ext_ssram_lane2_module;


architecture europa of ext_ssram_lane2_module is
              signal d1_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
              signal d2_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
              signal internal_q3 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 524287 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, clk) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;
    VARIABLE rd_address_internal : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    VARIABLE d1_rdaddress : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    VARIABLE d2_rdaddress : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "ext_ssram_lane2.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 524288) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rd_address_internal)));
      
			 IF clk'event AND clk = '1' AND rdclken = '1' THEN
                            rd_address_internal := d2_rdaddress;
                            d2_rdaddress := d1_rdaddress;
                            d1_rdaddress := rdaddress;

                         END IF;
                        


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity ext_ssram_lane2_module is 
--        port (
--              
--                 signal clk : IN STD_LOGIC;
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal reset_n : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity ext_ssram_lane2_module;
--
--
--architecture europa of ext_ssram_lane2_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal rdclock : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal d1_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--                signal d2_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--                signal internal_q3 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 524287 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--
--begin
--
--  process (clk, reset_n)
--  begin
--    if reset_n = '0' then
--      read_address <= std_logic_vector'("0000000000000000000");
--      read_address <= std_logic_vector'("0000000000000000000");
--    elsif clk'event and clk = '1' then
--      if std_logic'(rdclken) = '1' then 
--        read_address <= rdaddress;
--      end if;
--    end if;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "ext_ssram_lane2.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "REGISTERED",
--      lpm_rdaddress_control => "REGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 19,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q3,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            rdclock => clk,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q3;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library std;
use std.textio.all;

entity ext_ssram_lane3_module is 
        port (
              -- inputs:
                 signal clk : IN STD_LOGIC;
                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                 signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal rdclken : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;
                 signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal wrclock : IN STD_LOGIC;
                 signal wren : IN STD_LOGIC;

              -- outputs:
                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
              );
end entity ext_ssram_lane3_module;


architecture europa of ext_ssram_lane3_module is
              signal d1_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
              signal d2_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
              signal internal_q4 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
              TYPE mem_array is ARRAY( 524287 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
              signal memory_has_been_read :  STD_LOGIC;
              signal read_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);

      
FUNCTION convert_string_to_number(string_to_convert : STRING;
      final_char_index : NATURAL := 0)
RETURN NATURAL IS
   VARIABLE result: NATURAL := 0;
   VARIABLE current_index : NATURAL := 1;
   VARIABLE the_char : CHARACTER;

   BEGIN
      IF final_char_index = 0 THEN
         result := 0;
	 ELSE
         WHILE current_index <= final_char_index LOOP
            the_char := string_to_convert(current_index);
            IF    '0' <= the_char AND the_char <= '9' THEN
               result := result * 16 + character'pos(the_char) - character'pos('0');
            ELSIF 'A' <= the_char AND the_char <= 'F' THEN
               result := result * 16 + character'pos(the_char) - character'pos('A') + 10;
            ELSIF 'a' <= the_char AND the_char <= 'f' THEN
               result := result * 16 + character'pos(the_char) - character'pos('a') + 10;
            ELSE
               report "Ack, a formatting error!";
            END IF;
            current_index := current_index + 1;
         END LOOP;
      END IF; 
   RETURN result;
END convert_string_to_number;

 FUNCTION convert_string_to_std_logic(value : STRING; num_chars : INTEGER; mem_width_bits : INTEGER)
 RETURN STD_LOGIC_VECTOR is			   
     VARIABLE conv_string: std_logic_vector((mem_width_bits + 4)-1 downto 0);
     VARIABLE result : std_logic_vector((mem_width_bits -1) downto 0);
     VARIABLE curr_char : integer;
              
     BEGIN
     result := (others => '0');
     conv_string := (others => '0');
     
          FOR I IN 1 TO num_chars LOOP
	     curr_char := num_chars - (I-1);

             CASE value(I) IS
               WHEN '0' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0000";
               WHEN '1' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0001";
               WHEN '2' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0010";
               WHEN '3' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0011";
               WHEN '4' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0100";
               WHEN '5' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0101";
               WHEN '6' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0110";
               WHEN '7' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "0111";
               WHEN '8' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1000";
               WHEN '9' =>  conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1001";
               WHEN 'A' | 'a' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1010";
               WHEN 'B' | 'b' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1011";
               WHEN 'C' | 'c' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1100";
               WHEN 'D' | 'd' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1101";
               WHEN 'E' | 'e' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1110";
               WHEN 'F' | 'f' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "1111";
               WHEN 'X' | 'x' => conv_string((4*curr_char)-1  DOWNTO 4*(curr_char-1)) := "XXXX";
               WHEN ' ' => EXIT;
               WHEN HT  => exit;
               WHEN others =>
                  ASSERT False
                  REPORT "function From_Hex: string """ & value & """ contains non-hex character"
                       severity Error;
                  EXIT;
               END case;
            END loop;

          -- convert back to normal bit size
          result(mem_width_bits - 1 downto 0) := conv_string(mem_width_bits - 1 downto 0);

          RETURN result;
        END convert_string_to_std_logic;



begin
   process (wrclock, clk) -- MG
    VARIABLE data_line : LINE;
    VARIABLE the_character_from_data_line : CHARACTER;
    VARIABLE b_munging_address : BOOLEAN := FALSE;
    VARIABLE converted_number : NATURAL := 0;
    VARIABLE found_string_array : STRING(1 TO 128);
    VARIABLE string_index : NATURAL := 0;
    VARIABLE line_length : NATURAL := 0;
    VARIABLE b_convert : BOOLEAN := FALSE;
    VARIABLE b_found_new_val : BOOLEAN := FALSE;
    VARIABLE load_address : NATURAL := 0;
    VARIABLE mem_index : NATURAL := 0;
    VARIABLE mem_init : BOOLEAN := FALSE;
    VARIABLE rd_address_internal : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    VARIABLE d1_rdaddress : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    VARIABLE d2_rdaddress : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');

    VARIABLE wr_address_internal : STD_LOGIC_VECTOR (18 DOWNTO 0) := (others => '0');
    FILE memory_contents_file : TEXT OPEN read_mode IS "ext_ssram_lane3.dat";  
    variable Marc_Gaucherons_Memory_Variable : mem_array; -- MG
    
    begin
   -- need an initialization process
   -- this process initializes the whole memory array from a named file by copying the
   -- contents of the *.dat file to the memory array.

   -- find the @<address> thingy to load the memory from this point 
IF(NOT mem_init) THEN
   WHILE NOT(endfile(memory_contents_file)) LOOP

      readline(memory_contents_file, data_line);
      line_length := data_line'LENGTH;


      WHILE line_length > 0 LOOP
         read(data_line, the_character_from_data_line);

	       -- check for the @ character indicating a new address wad
 	       -- if not found, we're either still reading the new address _or_loading data
         IF '@' = the_character_from_data_line AND NOT b_munging_address THEN
  	    b_munging_address := TRUE;
            b_found_new_val := TRUE; 
	    -- get the rest of characters before white space and then convert them
	    -- to a number
	 ELSE 

            IF (' ' = the_character_from_data_line AND b_found_new_val) 
		OR (line_length = 1) THEN
               b_convert := TRUE;
	    END IF;

            IF NOT(' ' = the_character_from_data_line) THEN
               string_index := string_index + 1;
               found_string_array(string_index) := the_character_from_data_line;
--               IF NOT(b_munging_address) THEN
--                 dat_string_array(string_index) := the_character_from_data_line;
--               END IF;
	       b_found_new_val := TRUE;
            END IF;
	 END IF;

     IF b_convert THEN

       IF b_munging_address THEN
          converted_number := convert_string_to_number(found_string_array, string_index);    
          load_address := converted_number;
          mem_index := load_address;
--          mem_index := load_address / 1;
          b_munging_address := FALSE;
       ELSE
	  IF (mem_index < 524288) THEN
	    Marc_Gaucherons_Memory_Variable(mem_index) := convert_string_to_std_logic(found_string_array, string_index, 8);
            mem_index := mem_index + 1;
          END IF;
       END IF; 
       b_convert := FALSE;
       b_found_new_val := FALSE;
       string_index := 0;
    END IF;
    line_length := line_length - 1; 
    END LOOP;

END LOOP;
-- get the first _real_ block of data, sized to our memory width
-- and keep on loading.
  mem_init := TRUE;
END IF;
-- END OF READMEM



      -- Write data
      if wrclock'event and wrclock = '1' then
        wr_address_internal := wraddress;
        if wren = '1' then 
          Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(wr_address_internal))) := data;
        end if;
      end if;

      -- read data
      q <= Marc_Gaucherons_Memory_Variable(CONV_INTEGER(UNSIGNED(rd_address_internal)));
      
			 IF clk'event AND clk = '1' AND rdclken = '1' THEN
                            rd_address_internal := d2_rdaddress;
                            d2_rdaddress := d1_rdaddress;
                            d1_rdaddress := rdaddress;

                         END IF;
                        


    end process;
end europa;

--synthesis translate_on


--synthesis read_comments_as_HDL on
--library altera;
--use altera.altera_europa_support_lib.all;
--
--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;
--
--library std;
--use std.textio.all;
--
--entity ext_ssram_lane3_module is 
--        port (
--              
--                 signal clk : IN STD_LOGIC;
--                 signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--                 signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--                 signal rdclken : IN STD_LOGIC;
--                 signal reset_n : IN STD_LOGIC;
--                 signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--                 signal wrclock : IN STD_LOGIC;
--                 signal wren : IN STD_LOGIC;
--
--              
--                 signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
--              );
--end entity ext_ssram_lane3_module;
--
--
--architecture europa of ext_ssram_lane3_module is
--  component lpm_ram_dp is
--GENERIC (
--      lpm_file : STRING;
--        lpm_hint : STRING;
--        lpm_indata : STRING;
--        lpm_outdata : STRING;
--        lpm_rdaddress_control : STRING;
--        lpm_width : NATURAL;
--        lpm_widthad : NATURAL;
--        lpm_wraddress_control : STRING;
--        suppress_memory_conversion_warnings : STRING
--      );
--    PORT (
--    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--        signal wren : IN STD_LOGIC;
--        signal rdclock : IN STD_LOGIC;
--        signal wrclock : IN STD_LOGIC;
--        signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
--        signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
--        signal rdclken : IN STD_LOGIC
--      );
--  end component lpm_ram_dp;
--                signal d1_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--                signal d2_rdaddress :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--                signal internal_q4 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
--                TYPE mem_array is ARRAY( 524287 DOWNTO 0) of STD_LOGIC_VECTOR(7 DOWNTO 0);
--                signal memory_has_been_read :  STD_LOGIC;
--                signal read_address :  STD_LOGIC_VECTOR (18 DOWNTO 0);
--
--begin
--
--  process (clk, reset_n)
--  begin
--    if reset_n = '0' then
--      read_address <= std_logic_vector'("0000000000000000000");
--      read_address <= std_logic_vector'("0000000000000000000");
--    elsif clk'event and clk = '1' then
--      if std_logic'(rdclken) = '1' then 
--        read_address <= rdaddress;
--      end if;
--    end if;
--
--  end process;
--
--  lpm_ram_dp_component : lpm_ram_dp
--    generic map(
--      lpm_file => "ext_ssram_lane3.mif",
--      lpm_hint => "USE_EAB=ON",
--      lpm_indata => "REGISTERED",
--      lpm_outdata => "REGISTERED",
--      lpm_rdaddress_control => "REGISTERED",
--      lpm_width => 8,
--      lpm_widthad => 19,
--      lpm_wraddress_control => "REGISTERED",
--      suppress_memory_conversion_warnings => "ON"
--    )
--    port map(
--            data => data,
--            q => internal_q4,
--            rdaddress => read_address,
--            rdclken => rdclken,
--            rdclock => clk,
--            wraddress => wraddress,
--            wrclock => wrclock,
--            wren => wren
--    );
--
--  
--  q <= internal_q4;
--end europa;
--
--synthesis read_comments_as_HDL off


-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 



-- turn off superfluous VHDL processor warnings 
-- altera message_level Level1 
-- altera message_off 10034 10035 10036 10037 10230 10240 10030 

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ext_ssram is 
        port (
              -- inputs:
                 signal address : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                 signal adsc_n : IN STD_LOGIC;
                 signal bw_n : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                 signal bwe_n : IN STD_LOGIC;
                 signal chipenable1_n : IN STD_LOGIC;
                 signal clk : IN STD_LOGIC;
                 signal outputenable_n : IN STD_LOGIC;
                 signal reset_n : IN STD_LOGIC;

              -- outputs:
                 signal data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0)
              );
end entity ext_ssram;


architecture europa of ext_ssram is
--synthesis translate_off
component ext_ssram_lane0_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ext_ssram_lane0_module;

component ext_ssram_lane1_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ext_ssram_lane1_module;

component ext_ssram_lane2_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ext_ssram_lane2_module;

component ext_ssram_lane3_module is 
           port (
                 -- inputs:
                    signal clk : IN STD_LOGIC;
                    signal data : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal rdaddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal rdclken : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal wraddress : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal wrclock : IN STD_LOGIC;
                    signal wren : IN STD_LOGIC;

                 -- outputs:
                    signal q : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ext_ssram_lane3_module;

--synthesis translate_on
                signal data_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal data_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal data_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal data_3 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal logic_vector_gasket :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal module_input20 :  STD_LOGIC;
                signal module_input21 :  STD_LOGIC;
                signal module_input22 :  STD_LOGIC;
                signal module_input23 :  STD_LOGIC;
                signal module_input24 :  STD_LOGIC;
                signal module_input25 :  STD_LOGIC;
                signal module_input26 :  STD_LOGIC;
                signal module_input27 :  STD_LOGIC;
                signal q_0 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal q_1 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal q_2 :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal q_3 :  STD_LOGIC_VECTOR (7 DOWNTO 0);

begin

  --s1, which is an e_ptf_slave
--synthesis translate_off
    logic_vector_gasket <= data;
    data_0 <= logic_vector_gasket(7 DOWNTO 0);
    --ext_ssram_lane0, which is an e_ram
    ext_ssram_lane0 : ext_ssram_lane0_module
      port map(
        q => q_0,
        clk => clk,
        data => data_0,
        rdaddress => address,
        rdclken => module_input20,
        reset_n => reset_n,
        wraddress => address,
        wrclock => clk,
        wren => module_input21
      );

    module_input20 <= std_logic'('1');
    module_input21 <= (NOT chipenable1_n AND NOT bwe_n) AND NOT bw_n(0);

    data_1 <= logic_vector_gasket(15 DOWNTO 8);
    --ext_ssram_lane1, which is an e_ram
    ext_ssram_lane1 : ext_ssram_lane1_module
      port map(
        q => q_1,
        clk => clk,
        data => data_1,
        rdaddress => address,
        rdclken => module_input22,
        reset_n => reset_n,
        wraddress => address,
        wrclock => clk,
        wren => module_input23
      );

    module_input22 <= std_logic'('1');
    module_input23 <= (NOT chipenable1_n AND NOT bwe_n) AND NOT bw_n(1);

    data_2 <= logic_vector_gasket(23 DOWNTO 16);
    --ext_ssram_lane2, which is an e_ram
    ext_ssram_lane2 : ext_ssram_lane2_module
      port map(
        q => q_2,
        clk => clk,
        data => data_2,
        rdaddress => address,
        rdclken => module_input24,
        reset_n => reset_n,
        wraddress => address,
        wrclock => clk,
        wren => module_input25
      );

    module_input24 <= std_logic'('1');
    module_input25 <= (NOT chipenable1_n AND NOT bwe_n) AND NOT bw_n(2);

    data_3 <= logic_vector_gasket(31 DOWNTO 24);
    --ext_ssram_lane3, which is an e_ram
    ext_ssram_lane3 : ext_ssram_lane3_module
      port map(
        q => q_3,
        clk => clk,
        data => data_3,
        rdaddress => address,
        rdclken => module_input26,
        reset_n => reset_n,
        wraddress => address,
        wrclock => clk,
        wren => module_input27
      );

    module_input26 <= std_logic'('1');
    module_input27 <= (NOT chipenable1_n AND NOT bwe_n) AND NOT bw_n(3);

    data <= A_WE_StdLogicVector((std_logic'(((NOT chipenable1_n AND NOT outputenable_n))) = '1'), (q_3 & q_2 & q_1 & q_0), A_REP(std_logic'('Z'), 32));
--synthesis translate_on

end europa;


--synthesis translate_off

library altera;
use altera.altera_europa_support_lib.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your libraries here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>

entity test_bench is 
end entity test_bench;


architecture europa of test_bench is
component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc is 
           port (
                 -- 1) global signals:
                    signal clk : IN STD_LOGIC;
                    signal clk_to_tse_pll : IN STD_LOGIC;
                    signal pll_c0_out : OUT STD_LOGIC;
                    signal pll_c1_out : OUT STD_LOGIC;
                    signal pll_c2_out : OUT STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;
                    signal tse_pll_c0_out : OUT STD_LOGIC;

                 -- the_button_pio
                    signal in_port_to_the_button_pio : IN STD_LOGIC_VECTOR (3 DOWNTO 0);

                 -- the_cpu
                    signal jtag_debug_offchip_trace_clk_from_the_cpu : OUT STD_LOGIC;
                    signal jtag_debug_offchip_trace_data_from_the_cpu : OUT STD_LOGIC_VECTOR (17 DOWNTO 0);
                    signal jtag_debug_trigout_from_the_cpu : OUT STD_LOGIC;

                 -- the_ddr_sdram_0
                    signal clk_to_sdram_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                    signal clk_to_sdram_n_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                    signal ddr_a_from_the_ddr_sdram_0 : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
                    signal ddr_ba_from_the_ddr_sdram_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ddr_cas_n_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                    signal ddr_cke_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                    signal ddr_cs_n_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                    signal ddr_dm_from_the_ddr_sdram_0 : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ddr_dq_to_and_from_the_ddr_sdram_0 : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
                    signal ddr_dqs_to_and_from_the_ddr_sdram_0 : INOUT STD_LOGIC_VECTOR (1 DOWNTO 0);
                    signal ddr_ras_n_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                    signal ddr_we_n_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                    signal dqs_delay_ctrl_to_the_ddr_sdram_0 : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
                    signal dqsupdate_to_the_ddr_sdram_0 : IN STD_LOGIC;
                    signal stratix_dll_control_from_the_ddr_sdram_0 : OUT STD_LOGIC;
                    signal write_clk_to_the_ddr_sdram_0 : IN STD_LOGIC;

                 -- the_ext_flash_enet_bus_avalon_slave
                    signal ext_flash_enet_bus_address : OUT STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal ext_flash_enet_bus_data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal read_n_to_the_ext_flash : OUT STD_LOGIC;
                    signal select_n_to_the_ext_flash : OUT STD_LOGIC;
                    signal write_n_to_the_ext_flash : OUT STD_LOGIC;

                 -- the_ext_ssram_bus_avalon_slave
                    signal adsc_n_to_the_ext_ssram : OUT STD_LOGIC;
                    signal bw_n_to_the_ext_ssram : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal bwe_n_to_the_ext_ssram : OUT STD_LOGIC;
                    signal chipenable1_n_to_the_ext_ssram : OUT STD_LOGIC;
                    signal ext_ssram_bus_address : OUT STD_LOGIC_VECTOR (20 DOWNTO 0);
                    signal ext_ssram_bus_data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
                    signal outputenable_n_to_the_ext_ssram : OUT STD_LOGIC;

                 -- the_lcd_display
                    signal LCD_E_from_the_lcd_display : OUT STD_LOGIC;
                    signal LCD_RS_from_the_lcd_display : OUT STD_LOGIC;
                    signal LCD_RW_from_the_lcd_display : OUT STD_LOGIC;
                    signal LCD_data_to_and_from_the_lcd_display : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_led_pio
                    signal out_port_from_the_led_pio : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);

                 -- the_reconfig_request_pio
                    signal bidir_port_to_and_from_the_reconfig_request_pio : INOUT STD_LOGIC;

                 -- the_seven_seg_pio
                    signal out_port_from_the_seven_seg_pio : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);

                 -- the_tse_mac
                    signal ena_10_from_the_tse_mac : OUT STD_LOGIC;
                    signal eth_mode_from_the_tse_mac : OUT STD_LOGIC;
                    signal gm_rx_d_to_the_tse_mac : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_rx_dv_to_the_tse_mac : IN STD_LOGIC;
                    signal gm_rx_err_to_the_tse_mac : IN STD_LOGIC;
                    signal gm_tx_d_from_the_tse_mac : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_tx_en_from_the_tse_mac : OUT STD_LOGIC;
                    signal gm_tx_err_from_the_tse_mac : OUT STD_LOGIC;
                    signal m_rx_col_to_the_tse_mac : IN STD_LOGIC;
                    signal m_rx_crs_to_the_tse_mac : IN STD_LOGIC;
                    signal m_rx_d_to_the_tse_mac : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_rx_en_to_the_tse_mac : IN STD_LOGIC;
                    signal m_rx_err_to_the_tse_mac : IN STD_LOGIC;
                    signal m_tx_d_from_the_tse_mac : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_tx_en_from_the_tse_mac : OUT STD_LOGIC;
                    signal m_tx_err_from_the_tse_mac : OUT STD_LOGIC;
                    signal mdc_from_the_tse_mac : OUT STD_LOGIC;
                    signal mdio_in_to_the_tse_mac : IN STD_LOGIC;
                    signal mdio_oen_from_the_tse_mac : OUT STD_LOGIC;
                    signal mdio_out_from_the_tse_mac : OUT STD_LOGIC;
                    signal rx_clk_to_the_tse_mac : IN STD_LOGIC;
                    signal set_1000_to_the_tse_mac : IN STD_LOGIC;
                    signal set_10_to_the_tse_mac : IN STD_LOGIC;
                    signal tx_clk_to_the_tse_mac : IN STD_LOGIC;

                 -- the_uart1
                    signal rxd_to_the_uart1 : IN STD_LOGIC;
                    signal txd_from_the_uart1 : OUT STD_LOGIC
                 );
end component NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc;

component ext_flash is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (23 DOWNTO 0);
                    signal read_n : IN STD_LOGIC;
                    signal select_n : IN STD_LOGIC;
                    signal write_n : IN STD_LOGIC;

                 -- outputs:
                    signal data : INOUT STD_LOGIC_VECTOR (7 DOWNTO 0)
                 );
end component ext_flash;

component ext_ssram is 
           port (
                 -- inputs:
                    signal address : IN STD_LOGIC_VECTOR (18 DOWNTO 0);
                    signal adsc_n : IN STD_LOGIC;
                    signal bw_n : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal bwe_n : IN STD_LOGIC;
                    signal chipenable1_n : IN STD_LOGIC;
                    signal clk : IN STD_LOGIC;
                    signal outputenable_n : IN STD_LOGIC;
                    signal reset_n : IN STD_LOGIC;

                 -- outputs:
                    signal data : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0)
                 );
end component ext_ssram;

component tse_mac_loopback is 
           port (
                 -- inputs:
                    signal gm_tx_d : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_tx_en : IN STD_LOGIC;
                    signal gm_tx_err : IN STD_LOGIC;
                    signal m_tx_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_tx_en : IN STD_LOGIC;
                    signal m_tx_err : IN STD_LOGIC;

                 -- outputs:
                    signal gm_rx_d : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
                    signal gm_rx_dv : OUT STD_LOGIC;
                    signal gm_rx_err : OUT STD_LOGIC;
                    signal m_rx_col : OUT STD_LOGIC;
                    signal m_rx_crs : OUT STD_LOGIC;
                    signal m_rx_d : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
                    signal m_rx_en : OUT STD_LOGIC;
                    signal m_rx_err : OUT STD_LOGIC;
                    signal rx_clk : OUT STD_LOGIC;
                    signal set_10 : OUT STD_LOGIC;
                    signal set_1000 : OUT STD_LOGIC;
                    signal tx_clk : OUT STD_LOGIC
                 );
end component tse_mac_loopback;

                signal LCD_E_from_the_lcd_display :  STD_LOGIC;
                signal LCD_RS_from_the_lcd_display :  STD_LOGIC;
                signal LCD_RW_from_the_lcd_display :  STD_LOGIC;
                signal LCD_data_to_and_from_the_lcd_display :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_0_out_endofpacket :  STD_LOGIC;
                signal NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_clock_1_out_endofpacket :  STD_LOGIC;
                signal adsc_n_to_the_ext_ssram :  STD_LOGIC;
                signal bidir_port_to_and_from_the_reconfig_request_pio :  STD_LOGIC;
                signal bw_n_to_the_ext_ssram :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal bwe_n_to_the_ext_ssram :  STD_LOGIC;
                signal chipenable1_n_to_the_ext_ssram :  STD_LOGIC;
                signal clk :  STD_LOGIC;
                signal clk_to_sdram_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal clk_to_sdram_n_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal clk_to_tse_pll :  STD_LOGIC;
                signal cpu_custom_instruction_master_combo_a :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_b :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_c :  STD_LOGIC_VECTOR (4 DOWNTO 0);
                signal cpu_custom_instruction_master_combo_readra :  STD_LOGIC;
                signal cpu_custom_instruction_master_combo_readrb :  STD_LOGIC;
                signal cpu_custom_instruction_master_combo_status :  STD_LOGIC;
                signal cpu_custom_instruction_master_combo_writerc :  STD_LOGIC;
                signal ddr_a_from_the_ddr_sdram_0 :  STD_LOGIC_VECTOR (12 DOWNTO 0);
                signal ddr_ba_from_the_ddr_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ddr_cas_n_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal ddr_cke_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal ddr_cs_n_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal ddr_dm_from_the_ddr_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ddr_dq_to_and_from_the_ddr_sdram_0 :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal ddr_dqs_to_and_from_the_ddr_sdram_0 :  STD_LOGIC_VECTOR (1 DOWNTO 0);
                signal ddr_ras_n_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal ddr_we_n_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal dqs_delay_ctrl_to_the_ddr_sdram_0 :  STD_LOGIC_VECTOR (5 DOWNTO 0);
                signal dqsupdate_to_the_ddr_sdram_0 :  STD_LOGIC;
                signal ena_10_from_the_tse_mac :  STD_LOGIC;
                signal eth_mode_from_the_tse_mac :  STD_LOGIC;
                signal ext_flash_enet_bus_address :  STD_LOGIC_VECTOR (23 DOWNTO 0);
                signal ext_flash_enet_bus_data :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal ext_ssram_bus_address :  STD_LOGIC_VECTOR (20 DOWNTO 0);
                signal ext_ssram_bus_data :  STD_LOGIC_VECTOR (31 DOWNTO 0);
                signal gm_rx_d_to_the_tse_mac :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gm_rx_dv_to_the_tse_mac :  STD_LOGIC;
                signal gm_rx_err_to_the_tse_mac :  STD_LOGIC;
                signal gm_tx_d_from_the_tse_mac :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal gm_tx_en_from_the_tse_mac :  STD_LOGIC;
                signal gm_tx_err_from_the_tse_mac :  STD_LOGIC;
                signal in_port_to_the_button_pio :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal jtag_debug_offchip_trace_clk_from_the_cpu :  STD_LOGIC;
                signal jtag_debug_offchip_trace_data_from_the_cpu :  STD_LOGIC_VECTOR (17 DOWNTO 0);
                signal jtag_debug_trigout_from_the_cpu :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_dataavailable_from_sa :  STD_LOGIC;
                signal jtag_uart_avalon_jtag_slave_readyfordata_from_sa :  STD_LOGIC;
                signal m_rx_col_to_the_tse_mac :  STD_LOGIC;
                signal m_rx_crs_to_the_tse_mac :  STD_LOGIC;
                signal m_rx_d_to_the_tse_mac :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal m_rx_en_to_the_tse_mac :  STD_LOGIC;
                signal m_rx_err_to_the_tse_mac :  STD_LOGIC;
                signal m_tx_d_from_the_tse_mac :  STD_LOGIC_VECTOR (3 DOWNTO 0);
                signal m_tx_en_from_the_tse_mac :  STD_LOGIC;
                signal m_tx_err_from_the_tse_mac :  STD_LOGIC;
                signal mdc_from_the_tse_mac :  STD_LOGIC;
                signal mdio_in_to_the_tse_mac :  STD_LOGIC;
                signal mdio_oen_from_the_tse_mac :  STD_LOGIC;
                signal mdio_out_from_the_tse_mac :  STD_LOGIC;
                signal module_input28 :  STD_LOGIC_VECTOR (18 DOWNTO 0);
                signal out_port_from_the_led_pio :  STD_LOGIC_VECTOR (7 DOWNTO 0);
                signal out_port_from_the_seven_seg_pio :  STD_LOGIC_VECTOR (15 DOWNTO 0);
                signal outputenable_n_to_the_ext_ssram :  STD_LOGIC;
                signal pipeline_bridge_s1_endofpacket_from_sa :  STD_LOGIC;
                signal pll_c0_out :  STD_LOGIC;
                signal pll_c1_out :  STD_LOGIC;
                signal pll_c2_out :  STD_LOGIC;
                signal read_n_to_the_ext_flash :  STD_LOGIC;
                signal reset_n :  STD_LOGIC;
                signal rx_clk_to_the_tse_mac :  STD_LOGIC;
                signal rxd_to_the_uart1 :  STD_LOGIC;
                signal select_n_to_the_ext_flash :  STD_LOGIC;
                signal set_1000_to_the_tse_mac :  STD_LOGIC;
                signal set_10_to_the_tse_mac :  STD_LOGIC;
                signal stratix_dll_control_from_the_ddr_sdram_0 :  STD_LOGIC;
                signal tse_pll_c0_out :  STD_LOGIC;
                signal tx_clk_to_the_tse_mac :  STD_LOGIC;
                signal txd_from_the_uart1 :  STD_LOGIC;
                signal uart1_s1_dataavailable_from_sa :  STD_LOGIC;
                signal uart1_s1_readyfordata_from_sa :  STD_LOGIC;
                signal write_clk_to_the_ddr_sdram_0 :  STD_LOGIC;
                signal write_n_to_the_ext_flash :  STD_LOGIC;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add your component and signal declaration here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


begin

  --Set us up the Dut
  DUT : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc
    port map(
      LCD_E_from_the_lcd_display => LCD_E_from_the_lcd_display,
      LCD_RS_from_the_lcd_display => LCD_RS_from_the_lcd_display,
      LCD_RW_from_the_lcd_display => LCD_RW_from_the_lcd_display,
      LCD_data_to_and_from_the_lcd_display => LCD_data_to_and_from_the_lcd_display,
      adsc_n_to_the_ext_ssram => adsc_n_to_the_ext_ssram,
      bidir_port_to_and_from_the_reconfig_request_pio => bidir_port_to_and_from_the_reconfig_request_pio,
      bw_n_to_the_ext_ssram => bw_n_to_the_ext_ssram,
      bwe_n_to_the_ext_ssram => bwe_n_to_the_ext_ssram,
      chipenable1_n_to_the_ext_ssram => chipenable1_n_to_the_ext_ssram,
      clk_to_sdram_from_the_ddr_sdram_0 => clk_to_sdram_from_the_ddr_sdram_0,
      clk_to_sdram_n_from_the_ddr_sdram_0 => clk_to_sdram_n_from_the_ddr_sdram_0,
      ddr_a_from_the_ddr_sdram_0 => ddr_a_from_the_ddr_sdram_0,
      ddr_ba_from_the_ddr_sdram_0 => ddr_ba_from_the_ddr_sdram_0,
      ddr_cas_n_from_the_ddr_sdram_0 => ddr_cas_n_from_the_ddr_sdram_0,
      ddr_cke_from_the_ddr_sdram_0 => ddr_cke_from_the_ddr_sdram_0,
      ddr_cs_n_from_the_ddr_sdram_0 => ddr_cs_n_from_the_ddr_sdram_0,
      ddr_dm_from_the_ddr_sdram_0 => ddr_dm_from_the_ddr_sdram_0,
      ddr_dq_to_and_from_the_ddr_sdram_0 => ddr_dq_to_and_from_the_ddr_sdram_0,
      ddr_dqs_to_and_from_the_ddr_sdram_0 => ddr_dqs_to_and_from_the_ddr_sdram_0,
      ddr_ras_n_from_the_ddr_sdram_0 => ddr_ras_n_from_the_ddr_sdram_0,
      ddr_we_n_from_the_ddr_sdram_0 => ddr_we_n_from_the_ddr_sdram_0,
      ena_10_from_the_tse_mac => ena_10_from_the_tse_mac,
      eth_mode_from_the_tse_mac => eth_mode_from_the_tse_mac,
      ext_flash_enet_bus_address => ext_flash_enet_bus_address,
      ext_flash_enet_bus_data => ext_flash_enet_bus_data,
      ext_ssram_bus_address => ext_ssram_bus_address,
      ext_ssram_bus_data => ext_ssram_bus_data,
      gm_tx_d_from_the_tse_mac => gm_tx_d_from_the_tse_mac,
      gm_tx_en_from_the_tse_mac => gm_tx_en_from_the_tse_mac,
      gm_tx_err_from_the_tse_mac => gm_tx_err_from_the_tse_mac,
      jtag_debug_offchip_trace_clk_from_the_cpu => jtag_debug_offchip_trace_clk_from_the_cpu,
      jtag_debug_offchip_trace_data_from_the_cpu => jtag_debug_offchip_trace_data_from_the_cpu,
      jtag_debug_trigout_from_the_cpu => jtag_debug_trigout_from_the_cpu,
      m_tx_d_from_the_tse_mac => m_tx_d_from_the_tse_mac,
      m_tx_en_from_the_tse_mac => m_tx_en_from_the_tse_mac,
      m_tx_err_from_the_tse_mac => m_tx_err_from_the_tse_mac,
      mdc_from_the_tse_mac => mdc_from_the_tse_mac,
      mdio_oen_from_the_tse_mac => mdio_oen_from_the_tse_mac,
      mdio_out_from_the_tse_mac => mdio_out_from_the_tse_mac,
      out_port_from_the_led_pio => out_port_from_the_led_pio,
      out_port_from_the_seven_seg_pio => out_port_from_the_seven_seg_pio,
      outputenable_n_to_the_ext_ssram => outputenable_n_to_the_ext_ssram,
      pll_c0_out => pll_c0_out,
      pll_c1_out => pll_c1_out,
      pll_c2_out => pll_c2_out,
      read_n_to_the_ext_flash => read_n_to_the_ext_flash,
      select_n_to_the_ext_flash => select_n_to_the_ext_flash,
      stratix_dll_control_from_the_ddr_sdram_0 => stratix_dll_control_from_the_ddr_sdram_0,
      tse_pll_c0_out => tse_pll_c0_out,
      txd_from_the_uart1 => txd_from_the_uart1,
      write_n_to_the_ext_flash => write_n_to_the_ext_flash,
      clk => clk,
      clk_to_tse_pll => clk_to_tse_pll,
      dqs_delay_ctrl_to_the_ddr_sdram_0 => dqs_delay_ctrl_to_the_ddr_sdram_0,
      dqsupdate_to_the_ddr_sdram_0 => dqsupdate_to_the_ddr_sdram_0,
      gm_rx_d_to_the_tse_mac => gm_rx_d_to_the_tse_mac,
      gm_rx_dv_to_the_tse_mac => gm_rx_dv_to_the_tse_mac,
      gm_rx_err_to_the_tse_mac => gm_rx_err_to_the_tse_mac,
      in_port_to_the_button_pio => in_port_to_the_button_pio,
      m_rx_col_to_the_tse_mac => m_rx_col_to_the_tse_mac,
      m_rx_crs_to_the_tse_mac => m_rx_crs_to_the_tse_mac,
      m_rx_d_to_the_tse_mac => m_rx_d_to_the_tse_mac,
      m_rx_en_to_the_tse_mac => m_rx_en_to_the_tse_mac,
      m_rx_err_to_the_tse_mac => m_rx_err_to_the_tse_mac,
      mdio_in_to_the_tse_mac => mdio_in_to_the_tse_mac,
      reset_n => reset_n,
      rx_clk_to_the_tse_mac => rx_clk_to_the_tse_mac,
      rxd_to_the_uart1 => rxd_to_the_uart1,
      set_1000_to_the_tse_mac => set_1000_to_the_tse_mac,
      set_10_to_the_tse_mac => set_10_to_the_tse_mac,
      tx_clk_to_the_tse_mac => tx_clk_to_the_tse_mac,
      write_clk_to_the_ddr_sdram_0 => write_clk_to_the_ddr_sdram_0
    );


  --default value specified in MODULE button_pio ptf port section
  in_port_to_the_button_pio <= std_logic_vector'("1111");
  --the_ext_flash, which is an e_ptf_instance
  the_ext_flash : ext_flash
    port map(
      data => ext_flash_enet_bus_data,
      address => ext_flash_enet_bus_address,
      read_n => read_n_to_the_ext_flash,
      select_n => select_n_to_the_ext_flash,
      write_n => write_n_to_the_ext_flash
    );


  --the_ext_ssram, which is an e_ptf_instance
  the_ext_ssram : ext_ssram
    port map(
      data => ext_ssram_bus_data,
      address => module_input28,
      adsc_n => adsc_n_to_the_ext_ssram,
      bw_n => bw_n_to_the_ext_ssram,
      bwe_n => bwe_n_to_the_ext_ssram,
      chipenable1_n => chipenable1_n_to_the_ext_ssram,
      clk => pll_c0_out,
      outputenable_n => outputenable_n_to_the_ext_ssram,
      reset_n => reset_n
    );

  module_input28 <= ext_ssram_bus_address(20 DOWNTO 2);

  --the_tse_mac_loopback, which is an e_instance
  the_tse_mac_loopback : tse_mac_loopback
    port map(
      gm_rx_d => gm_rx_d_to_the_tse_mac,
      gm_rx_dv => gm_rx_dv_to_the_tse_mac,
      gm_rx_err => gm_rx_err_to_the_tse_mac,
      m_rx_col => m_rx_col_to_the_tse_mac,
      m_rx_crs => m_rx_crs_to_the_tse_mac,
      m_rx_d => m_rx_d_to_the_tse_mac,
      m_rx_en => m_rx_en_to_the_tse_mac,
      m_rx_err => m_rx_err_to_the_tse_mac,
      rx_clk => rx_clk_to_the_tse_mac,
      set_10 => set_10_to_the_tse_mac,
      set_1000 => set_1000_to_the_tse_mac,
      tx_clk => tx_clk_to_the_tse_mac,
      gm_tx_d => gm_tx_d_from_the_tse_mac,
      gm_tx_en => gm_tx_en_from_the_tse_mac,
      gm_tx_err => gm_tx_err_from_the_tse_mac,
      m_tx_d => m_tx_d_from_the_tse_mac,
      m_tx_en => m_tx_en_from_the_tse_mac,
      m_tx_err => m_tx_err_from_the_tse_mac
    );


  process
  begin
    clk <= '0';
    loop
       wait for 10 ns;
       clk <= not clk;
    end loop;
  end process;
  process
  begin
    clk_to_tse_pll <= '0';
    loop
       wait for 10 ns;
       clk_to_tse_pll <= not clk_to_tse_pll;
    end loop;
  end process;
  PROCESS
    BEGIN
       reset_n <= '0';
       wait for 200 ns;
       reset_n <= '1'; 
    WAIT;
  END PROCESS;


-- <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
--add additional architecture here
-- AND HERE WILL BE PRESERVED </ALTERA_NOTE>


end europa;



--synthesis translate_on
