  --Example instantiation for system 'NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc'
  NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc_inst : NiosII_stratixII_2s60_RoHS_TSE_SGDMA_sopc
    port map(
      LCD_E_from_the_lcd_display => LCD_E_from_the_lcd_display,
      LCD_RS_from_the_lcd_display => LCD_RS_from_the_lcd_display,
      LCD_RW_from_the_lcd_display => LCD_RW_from_the_lcd_display,
      LCD_data_to_and_from_the_lcd_display => LCD_data_to_and_from_the_lcd_display,
      adsc_n_to_the_ext_ssram => adsc_n_to_the_ext_ssram,
      bidir_port_to_and_from_the_reconfig_request_pio => bidir_port_to_and_from_the_reconfig_request_pio,
      bw_n_to_the_ext_ssram => bw_n_to_the_ext_ssram,
      bwe_n_to_the_ext_ssram => bwe_n_to_the_ext_ssram,
      chipenable1_n_to_the_ext_ssram => chipenable1_n_to_the_ext_ssram,
      clk_to_sdram_from_the_ddr_sdram_0 => clk_to_sdram_from_the_ddr_sdram_0,
      clk_to_sdram_n_from_the_ddr_sdram_0 => clk_to_sdram_n_from_the_ddr_sdram_0,
      ddr_a_from_the_ddr_sdram_0 => ddr_a_from_the_ddr_sdram_0,
      ddr_ba_from_the_ddr_sdram_0 => ddr_ba_from_the_ddr_sdram_0,
      ddr_cas_n_from_the_ddr_sdram_0 => ddr_cas_n_from_the_ddr_sdram_0,
      ddr_cke_from_the_ddr_sdram_0 => ddr_cke_from_the_ddr_sdram_0,
      ddr_cs_n_from_the_ddr_sdram_0 => ddr_cs_n_from_the_ddr_sdram_0,
      ddr_dm_from_the_ddr_sdram_0 => ddr_dm_from_the_ddr_sdram_0,
      ddr_dq_to_and_from_the_ddr_sdram_0 => ddr_dq_to_and_from_the_ddr_sdram_0,
      ddr_dqs_to_and_from_the_ddr_sdram_0 => ddr_dqs_to_and_from_the_ddr_sdram_0,
      ddr_ras_n_from_the_ddr_sdram_0 => ddr_ras_n_from_the_ddr_sdram_0,
      ddr_we_n_from_the_ddr_sdram_0 => ddr_we_n_from_the_ddr_sdram_0,
      ena_10_from_the_tse_mac => ena_10_from_the_tse_mac,
      eth_mode_from_the_tse_mac => eth_mode_from_the_tse_mac,
      ext_flash_enet_bus_address => ext_flash_enet_bus_address,
      ext_flash_enet_bus_data => ext_flash_enet_bus_data,
      ext_ssram_bus_address => ext_ssram_bus_address,
      ext_ssram_bus_data => ext_ssram_bus_data,
      gm_tx_d_from_the_tse_mac => gm_tx_d_from_the_tse_mac,
      gm_tx_en_from_the_tse_mac => gm_tx_en_from_the_tse_mac,
      gm_tx_err_from_the_tse_mac => gm_tx_err_from_the_tse_mac,
      jtag_debug_offchip_trace_clk_from_the_cpu => jtag_debug_offchip_trace_clk_from_the_cpu,
      jtag_debug_offchip_trace_data_from_the_cpu => jtag_debug_offchip_trace_data_from_the_cpu,
      jtag_debug_trigout_from_the_cpu => jtag_debug_trigout_from_the_cpu,
      m_tx_d_from_the_tse_mac => m_tx_d_from_the_tse_mac,
      m_tx_en_from_the_tse_mac => m_tx_en_from_the_tse_mac,
      m_tx_err_from_the_tse_mac => m_tx_err_from_the_tse_mac,
      mdc_from_the_tse_mac => mdc_from_the_tse_mac,
      mdio_oen_from_the_tse_mac => mdio_oen_from_the_tse_mac,
      mdio_out_from_the_tse_mac => mdio_out_from_the_tse_mac,
      out_port_from_the_led_pio => out_port_from_the_led_pio,
      out_port_from_the_seven_seg_pio => out_port_from_the_seven_seg_pio,
      outputenable_n_to_the_ext_ssram => outputenable_n_to_the_ext_ssram,
      pll_c0_out => pll_c0_out,
      pll_c1_out => pll_c1_out,
      pll_c2_out => pll_c2_out,
      read_n_to_the_ext_flash => read_n_to_the_ext_flash,
      select_n_to_the_ext_flash => select_n_to_the_ext_flash,
      stratix_dll_control_from_the_ddr_sdram_0 => stratix_dll_control_from_the_ddr_sdram_0,
      tse_pll_c0_out => tse_pll_c0_out,
      txd_from_the_uart1 => txd_from_the_uart1,
      write_n_to_the_ext_flash => write_n_to_the_ext_flash,
      clk => clk,
      clk_to_tse_pll => clk_to_tse_pll,
      dqs_delay_ctrl_to_the_ddr_sdram_0 => dqs_delay_ctrl_to_the_ddr_sdram_0,
      dqsupdate_to_the_ddr_sdram_0 => dqsupdate_to_the_ddr_sdram_0,
      gm_rx_d_to_the_tse_mac => gm_rx_d_to_the_tse_mac,
      gm_rx_dv_to_the_tse_mac => gm_rx_dv_to_the_tse_mac,
      gm_rx_err_to_the_tse_mac => gm_rx_err_to_the_tse_mac,
      in_port_to_the_button_pio => in_port_to_the_button_pio,
      m_rx_col_to_the_tse_mac => m_rx_col_to_the_tse_mac,
      m_rx_crs_to_the_tse_mac => m_rx_crs_to_the_tse_mac,
      m_rx_d_to_the_tse_mac => m_rx_d_to_the_tse_mac,
      m_rx_en_to_the_tse_mac => m_rx_en_to_the_tse_mac,
      m_rx_err_to_the_tse_mac => m_rx_err_to_the_tse_mac,
      mdio_in_to_the_tse_mac => mdio_in_to_the_tse_mac,
      reset_n => reset_n,
      rx_clk_to_the_tse_mac => rx_clk_to_the_tse_mac,
      rxd_to_the_uart1 => rxd_to_the_uart1,
      set_1000_to_the_tse_mac => set_1000_to_the_tse_mac,
      set_10_to_the_tse_mac => set_10_to_the_tse_mac,
      tx_clk_to_the_tse_mac => tx_clk_to_the_tse_mac,
      write_clk_to_the_ddr_sdram_0 => write_clk_to_the_ddr_sdram_0
    );


