��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ��p"���C��T�fX��k�+��)��6�'�3��$���)��2�+�
�#�7��Ib����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`lJ�g����BĬ������M?Ŋ�#��I^����b�,ozz-h3�D�r[k�j2�'���`�<g�k�K��q3ŭ�NĮ4�Y���F?O�vI�M�|�TZ]�!��s6����*[3���Y<�D&��cP�]�{�s2p��E�哦=��dG��UKR����#�^��J�T���Q��р{��\5x��'�@�_��?�� L�HQ+o�)����U��b�e��im�R-�6�Y�O�� o��;�"R�m^�w*��F���E�]NX��������z��#K���|{
��+��8ҁ�-桖��$]�����G�H$�]gvVw$9̳�N�Ӵ�!�r|�~�ZGU�1=�Qz=�T��@�nN3�{�����Go�l�X;�]���Պ���,��%1�Y�|�V�!H�<l�[8:4 ��{5�SQ�*٠�\��G� ¸�9�2'N?"�U���C4Sw�RxQR�dYP��HѿӅ+�Y4���w������x�A@�����р�Pw�W��W��6D�����bJL�!�}��2<��H�c���U�ˬ�>n���|��MWAD%��9�1�����"F�3x	�������Btd���5�Pj+��6u������ֆx��Wi޶�!��CX���J���G���s&��dM5���f3��"x� x
8Ǣ�Gö��?��TN��
�ܯٵ,J�h��v���/b���_���"�1e��24�P�sJJ�*.�̑a�B ���'�U#�]�1���W�� �3�j���I�~;�>��ǓB�Xb����Zf�@�\�P\�����ܨ��������vGHQ+�2�@�ƹ\�8���Y >�4	/DZ>�Q?��D硫���S��[�`ވ<���w`'�{����u�>Ѭ�Ķ�<eǒX���
t�5F�r�;���5#x�`�L��-Ni�!��	���i���蕐�;���oɜ7�u��b�!͐��q�I
nj�$��r��u��-ft��-74������B�����"��jD�_�ܣKpJ��_<�2cxT�[X�\�꘺�hn(t��cR�zI�-�B�zg�<hӔ�̓ȜǬZP��H1iΘ6���%��A7��=�C��]W��wN�ti��FXZ�
�EGGת�-F�|"�-�
�_fm]�^�va�ǰ>㷵��� yD�s�<���.p\�/;h7��:�K)���QBJ΢)D�xb�I
\�8sd� t��{�]z�R������!*����<@��s2�P����}��|�ס����l����"T�)����6}���7 �h	;dF��Ӹ	�MWrL�G ��߶�5���k���ꇅ-4�z��YT�C��!k�/>�� ��I�XI���d�7�·�ՉB�W�b*�6��e"�U�r�t�2���9�ZX�`gP�O*<}�1$re5K�]�[�f�vX�E���{�7FOj4*\�f��Q6��n�{>3�
~���fƿa��U��*\0_�OU�%���ņ�!�v�]��:͹A��r������Y��� *n��0�M�=Vk��1���![�,,��u�^����;�n��ٗV����z{�|-a�ĕ�@�R��v�3W���:�c���A��{0����J�(�ݨ�H���֯�l�m(@3)u�E?Nk]G��Cࢾ�k�\�ݕLW��ծ��>���w6��v��ڹ|�M�͊�Y��v\�����L���Ω����JW�`c���4��%�X�%�"qzcgN�� �}	k��5�()4I?�	�E�7��?�_�_�ɣ��Fi��72�Cj1۠���=�*��)i1��+\���s҆d�'A�iT��3nt�AZ��#j#KB���@k�7�H�D�s_�F8j�� ���`�|�!��mU�J(�ۼ�"�Vu�} #RK���S�	n�ydbZpY��0/ۇ��^��z�K�������*�Xי��lcJ�oΙ�{��`8�6��i�!���_},�?�"5���������v���8�xfHK�@Ě1�Ή.�Xz��G�]O�ݺ�[֨��*�z�嘭ε��9���!^`��}`[Lv$�#4�<@�ζ�g�dC{��ڌ+ 7��g<��!G}�؝7�7<�EA��۬+^���^�B��l�_��.�+'䃹{���t~XC���-!����ԏW���2+A���79��Di���o_��>|���,1*N��<�'(q���gbtߓ��:��46B��7����}l/b�-{�f&���K��Ȧ�b��6IZRN��Ĉ�򊭅@��4���%A¡�D��geJ��g����Y���z���u�K�T����$@-J@��5ʙ3G�D�$����O�����՞��_���s$0���>]��`�|D�:Zq~VҺ��DU Z�ُ�<�Q�)F-� ����5h�D�.nhB�TU�Pa�Q�2�A�H_
��
��[?b�8B�����:���-t�:)�,�胓�I��dUӰ�ŝnq�I�uNqռ� ��y����e��+K�� �3�D����R~���U"Tㆧg�X��Y�q�X�THm:ݲ7�f��� ��5�a�ؖ���촄G�W�#I��&^�Da+�C�$?!�������&��u4賀��oo��yߢ�#L�3�3���*�vy,\��7DMF����D�o������K�E���(c�sC�5?�߮� �9����*r�i���y�'\]%�h"B0�� }$.%+d:ʠm� ���.v����o�]`�`��T^cI_�z �Dc�SǮ5-�5��Sd�e�ԛ�n����Z{�����E���n�](����֑_o�R�xq��Pg_=�諪KH.��/��n��^�������
�{��x"P��q�;�^@h6g�l�ce�N�Zk��	�)���}s�fi�X�V�8i���̚��D%c��!p�7@	�f�J�I�Т�%	c���J�ɴ0�����־����u1������HA�"��:_]�%��n
���i-�A�����7�ղ![�/�b9���2J����`,.�{%6�#ݷ!D_� m�����Z��A�͑8�+w��a�m�Y����g� ����E�)Ʊㄱ�6`���3PgP=��*�����,�����샞��G�O^��y��@�%���4��-p�i8���z���'$��1{��C/5�1���$����=��*�����Tn[c�ލ�yy}]�v i�0fl�Ҍ��8*���
e �������b�b_��C�|��y�R�_Sg����Wǻ��KWd����.y���%U�B�'%k�6Py>�sS.�ⲣ�~��i'������&.��7�I)M��$`��C�6�	�G�|0���w�t���E�-����s�No!��v͠�ce�	��2Ŷ#3��Ig+��lO���I�j(�R7�b����"�O��2��-�A<��U��@��YC
GZ(�Ū�});�e��Er#���a^���s���~/���ü�NѸɭ�n���簑�O*.��,�w	$��H-�������b�Z�x�C�m��D軂�V���JR����`��E���HD��ǳt4��N�?Wٌ}�@WBچ�5�t�����3��¹|�
����_i'C�>��j'�U�ű�*����A����ǫ���='�%ӵ[��U�a�}����;�ҙ�g�NKk��Ǿ��;����Î����=Fd�ګ{��xĀoWM�l����x�#�,_��Ç,9�Q��)~���o�N������%`�k	��F�Gg@����"	�j� �M����}�oT��؊��R�^�`���0��:�Z������0,�z��
�7]/ѭv轛6���I::�&=K�B�=虮����"��X r�V�# P?�C�NӉ����GVtPvC1Wz�Rd5�OC�z]D�K�~VE��i˦2b9j|�BI�A��j�Tӱ}r/���$,+�̤^70QCY�Nq�!tc�qJ ���]� l%��<��>�����T����:���F�/	�\^��4�����C0��P�̧4S{���@4� �97�[duk^[3su�gx���]�Um&s�[�A��u��_���5r�@0��#����펈DJ�)bK�1��S��G�������p���̼=dw�@Je�nR��q+8ɕ�ո:)U0_�.� �5e�l����?�2�so������F�3&{mb��H$~$fE)F�2f.��/��H�� �cу.P3e�Q��w5�]�ÖS��T�[{8b^�)��؏���xL:�`���(�_��4�bS.k|sd���ċt��뻖\��P>��y¢.k��Za�ہ��Q ��vh�G���H��o	��t��2�B� $� ��y��v@0�ò��ݥ��따� ��{s�,�Ԭ+��X���6��%����j�*L����qٴ_��ի����ϒi�M��T��F�>pp%ń�w����T��Hm����mܶh�|�i 5��Q1n�,�Q�!l~�l�̢S·���?�;���Z=t��<���sRq��H�Gc:Ϛ��.p��0R�w��C2�9��c	�*] =RF'=�b�{���Vz&؈���L��Z�[�#��v�Z�%�
v�_�/�?�,h�jY%]�`[����A�A�����VZ�q�z�!��;��v�Ȓvf(]��v�$�sk�f�;�A%2�k��K��ƥ�duT�~��9���u3[�0Ym�M���=�H2Lz��8١�LO���B.���fQ�OT���O�?D�cb����D�x��3��Br[���I?��l��E�%�.�\��bFRKtߘC|���=]��x��������o:������vJ�;��!��S��J��w75�5o�{����W���.$!�#�	)��7|4�4���$��.	%�mک���W�������~@ϩ71��M��Ip� z�����{�/e�
{�?��7D>�W�C�<>k�7l����|ݻ�Z(�~���L�2K$X9�o)hH��.w��|�Y�ۘ�4�N^�g�����s^~&1L�a�hw�-1F�7�"�@m��+�w��S����[/؄�^�;R�S��XʶٽM����pD��,�}��¹�`E7���o��#'���7�˯wRS�Ϯ����f�D^ws��Q��@��hu?ѩɝ Ddm�&/��%�9N࣓H��B�+�������{�#O�+ؘ��
�AU`�-A�,k��j�ɤT������D*�o��1(;�Mϭ�X&
Y̝�]�t���������[���vڰd$q �`��F!"#���i�� =C���X'�Ƥ�}.JO����jG��z�>7��D��Ҽ`�k�����28 �����Ԣ��"�n�N������_IZR=�rP�gI;h�T�9dfHF+h�N�`qf�Èv�!z
=��n:A���9Z�*Nv�� Z���b���Js6���`�T?ܷX���!�j�k]����������՛ ��H���
�k�hu�������r�/!Yj�6q"��A��nk��AT�qH�&�"=$�֏*�g�X�.�\K=���s��%�,�U'��M@=��Rm#�W fm������ɐˡ:A zi.P؜fZV+�
M[��0��r���}���
���Yb[5�&:��C��F�M�L����0�l5���x���������&8Q`Z"KM�D5]�=2���h��� d�����������˕�H�7��w���nu�~��(�!���
f�ׂ&��|�\,_�7�� <0(wFfTm��<���YK��wR6`Ja�E�T��#�ڏ)qE�Z+�;���wzAFT�>�+U��Kµ���kQ+�Z����t�X�E�#5X�`9�C)9s_T,��/~��t)��ϩR�����g�X50��E��D���Y�G�� ��,�;ґ�?�QV~a��Oՠ�Ϛ7q��	�y�x����D|��˘c�"��:���jܢl��.׊<rɄz��i�K�#����G��t�ٛ�a�1t[w�^�b�	$}�i�.�"F�V�t�n���d���-���; �����LR�W�(s`כ��������/�(�U�եо��YNw��V�	'����W�ʬ�I$E������φ��	�%sw@�@�㫙<�;~�q�;�>W8���s�e2�����"d�p\�X�1�m�x�w���Ͷv�����:��<,�����o�Qy�{���K�mp��t��sw�8R�Y_����<p��������e���7CT�6�=����6�5?��e�k�<�Wf�qdb����1{N�M!�J�s�F�)���b�jw�����)c_�v���Om�6���H�5�3�qT�qh�䈩-�Y������o��F�`|+�w���*��Ԏi���9��Ü�%|�M_�Z���eI�N�:���w��;�iFUѰ�m�,����QH 
��]���2^j/�����@[W;z�~��d^��ț�y p��^7���Y�i8��ِ����{A�xAM��9�d@m!� }�A�˰%���x��b ����ݡ!�h 1��d*<s�2hq%��D�������pȅ��o>�����vօ�Z |1��H�f�U�>�)J߱��x�b�s�="'����E�*6.,�)�'���^��Ej��җ�}M�%z"�K�lX�U(�l^�{k���{c�۝&_�(���/$&����O��p!�A�$X��:/�vB��f���-��M�KV���	h�S����n�Bs�hlN�˷��FZ�$G0�$l�o���[���;�y�~��o���:\�'"Y_��ɗ.H1�.�&������ك�Z���Wؘ�ckS����zy �)�Ӽ0��9ԉ9�Ğ8&bQ���Q���fm[�R"3L!_(�!(�.��<}X�-i�~�4�u	���.c�qo��|�5��0�*�ї����$G��`-����/�mH]#�׸���Z�`#�jI��R�G�l��C��թa@W���f��@A
��r�ѷ��ʕ�Oә�v��wڣ|�ड़���g�R:@l��򵿛��~�͏*��b!��ߌ�\Y�{FAŵ�.��|��;�?'�vL��(�MN�y���X1�q�;v�3Nw��*|�5�;�;<��i������o��m�V0A(��_�@ �9�x��Ȉ��ݢd�HM������Ħ���Ɩ�
k���7���Dd�+�mY��|����y^  ��;���y	A@�����dM��1�5!Z\M�����z"h�xٛ{� %��_���!¶S^Z��x��^g�Rަ��GB ��=_7@/ �g%�%��I��pX�,p�ڬ9ǀḘ�ݔ�q��1ޣ��j��'ѫ��J��������m��k�jk�U���Վ=$k�8D��T;����]n�6�ٯ�U����ݞ��	�R��:	�o�ڟ��Bdh�5��ղkȑ�=_K�sE>��s�,��'���J8�r%��-��@<`�sK\�]��������	I�W�gO��M�Q��y]<c~Di��߸�5����F_��K���+���"DyV,C,
gH=h?��M�}䱒} � �^U6m5c�������8ʊlP�̘�E����j�%v~��a34�QyK
�eNUMo'��
�����F79!i
��+S��[.�-�D��^�,�ʩ�# r�M�MœZ��X�iY4`ţ; ą<JH3K]%�C�i��$j3U����W��%�ɢ��و��X>o��t�Q�1}�F�S��ϙ�-�m~\�n؊ �a���1�0�&���Qk/�<�R�΁d�L �Oݓh�-@ ���!#�]/M`0���6��;��߹<��%�gi(i�kxb5\�`���k�P�D䁠ZZ1U0}/���:7*���x���A_�� P��0o��Վ�z
��u�<�W�{�B��5�<ͻª�*�[�}��^'HːaA���'`!^�4QR��e���O��T�����@�[U�|Q��:1�&��!�|� #��FM8����a�6�/P<yi%�ջ�D)�nH��h�������UU`�a&�G!6O��%�~���� #VH�RB�#p�ƒ�\u�G���������Sg���*�,�D[��=�{:u;Q��,����Z�{^j�'�Q��
��-��?ь�o�KPZmGO��2�|���[�h���$���ׯA^�]���gq�Ɂ��?c
�@�4�4X".��W����j8�պ�$wK�x=QW�h$�3��ʋ��4zΠ�q��"?^IbG�����1�i���*f7u�����[���;F�B��Jw�������Z�����\�	�3ܑ99ӈ�^��Y���;J����_Ȃ�@+&`�ڑ\=�,2질�D�h��=�-�}�B�]5$�d�"�������J	\��r���^X\����u�!�EPsj ���=��[����������y	iH&pQ��\��U�S�v��]ƛV��\{)�j�Uf�D��g�DV�c����Sl��1^W��
}G�
�j~�O���4^�󯫙�M�<�H Lg��{ǋKb�^=�O,q�7k�6��Z�İV�.���g7�;W�
�	�:7��^�l�T�<�]C��x���A�Qw�'p�h�9d��,G�R!�4��4e'�`��I�����%Y�~P|�t������!u0��#�@!�T{NӇ��)�L.���M�X�Մwϓ)ygg�_J��� ߄V4N�]c���]���C����p�T���<6����M0�8�C�����z�����1��yY] ����TD;Ӵm��)5\y���� �-k�z֏h�Ci�$�@�����)���m��uY88`oφ��Q7��?�AI�ל���ߵ�R6��'|�?iɾ�
��OVl٭ф���E5T����yl�K���"ok�Ҹ�q qVs5���h!�(1O�4-�9�C]�5���x��b�|�[��ŏ,[mrW�[N.��P����b#K��a�:y70B���%�x��>>D�[W���d����_��k .�SVP���LvĞ��.��<Q>���%r3��[��&;]���vi��Xgg�-���T:R�ǂ�l�w�U��DJ�m��'��㗚�b���n*���v�W[ܬ�nAj�tZ��rJ�<4B�;��ut��:cm �O\�(����W޿&V�]P8��:ͅ��Եq��Ղ�YJYL�P0`!�����!���\c.i!iv!:}׳)JǭM�s�9��3J��I�,�7Q�o��5��J��/����\b��}�J>9g`��}g��/P��E���J+��b`
AO�q��/I��D�3m�+����d⒚���֝�������k@!���'��j�=�c�U؜L�џ/5hG0��l=f��'� ���߶K������C���=�����
�,P��j�%�~�[���RB]�p�+�g:�\ԁ/8�_�mkDsf�ԌACzY� I�,tdu�zsU�t��(7�C9Ģ�?Uj4�ةZWFש}� uv�C���|͵)␦��d�rO��������m�.�<p�*)G#�ݽ
$���6'�5L��X*{���TJrlD�� �X�gwJ>��r]75I����\���?sBz���[/6�)ֿݵ�ͣG���а�CP:�0y�>O�O͜����vy<�A'Mၤs
:�v�o�i���}b� �h�������z�}u(ħ����*K���fTNi��u�F���s1Ĕ�Җ�(R�u��r0l�X������2!ͅ�	$e
M>�k����ĜSf\A]�����I4��Ƽ�}�g��n7C��4]u2��㬉����o�0Ǒh̰T<�j���X.DY�$	`(ٚx�n0��Ҹ�W0X�.����?��!�s�;7Q�a��BO��W�j�;�(�J�� �?$��_�e�����b%Q�Y�^w����DX�_&�#jS��Ŏ�ܬ�O�<�+Ʈ�)��F�6n�G��I.��8���C�S�����A��4.AU�#.� ��J(�ذ5�4X�T00���S��H����ʱZ��r{_=��+j!�]�R��)S��]^	��3M9��5-��M�l�۹J��I�Ҿ��I����}�)�N4/|�2�`6q)�9��H��ư�T��y�T�_F���'`��/�-]"*0^N�U盛��[8`U�)E�tБ:��q,9?gY�ib�O9�ܩ	ּ��Y����+H=ϛ���K`[)A�N��R����Ѣ1>B^�ch��%�&�༁5����mN��,�Ph�t�a�A�U`�O��
6�Çs+����>c�S�\���0�]J}������x�O�^���2�̤]3 �z��/��L/���R��	&
)V4&�����UQ��ͧJ�{���JC��b(�fq|��%�	�b����̒�~�ॽ6��	�����t�&ކ����'��f�1>��)��a�cS�a��1c{����`����3�P`�{�!me6c�U۳5�3'�!y�yT��K���f/�/mj
`I��8�%�������i�E�6<�2��z�cW� i���7vCӠ6`�.:�5+բ�$I
gK��,��0��"E�r;�e��)����'�Xm���yE-K�I.ߣ�	r��̅�bϳ+m�a�f>e� �ͺr S����<�)�Ӛ�i��� �=������M��2@��F�c�1�FM9���a���С��7�q��r)����Vdlr�_���̲Ql?kF�zcG\GF��R�ɑ|�7�q�����N���X���^�U��Zj �@S�oB,�p�G�^.���fb�V��.Ŧ1{���u���N��2)