��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ��p"���C��T�fX��k�+��)��6�'�3��$���)��2�+�
�#�7��Ib����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�Ē\dEkU�n�]7K��	S���(}�,Ϳ-�n�U��;]րi���;$vdm�	�M����-[r��'Y�r*|�2{t��V �X�<M|�z��Z�۳�&F����~U�N�w��b�&?�@�V�Bm+Up���:�l��i/z4�YS�Pm���f�O��9�B��ػ�ɪ��g�(R�A�gBM�AB����kV�(�i|��!.�C1�^!��1P�i��$J��Y�Q��(��tԂ~-�XTW��?(�]�6�؁�X�@U���H��je�`	��j������/a�jqȏ��5BY ؏����?����MR\���L���k� 8`B��'}p���L]˃�h]A�����F�&�&3ا�i#�TZ�5��}8�ʏ}t�>�#���C�_��6ꏉ\m�M�vVy^���iH8�_�(�ĈC���Hߢ����% n�C��K�����D�ٴ+e�q�q���x��X�]}%��#�6=����+��3Y��lP��U��/�����%���& g7�c��4����?�W_�!3�k ��紴���x��T��ۙ^�k���h�ؘ�B6�T՜�֔� ���N�'P�Pb��B��(	�;=�^���~L3R^�Y����C�?M�_���H�*��\�^z%��ٗ��/����`�Ko䓿��E����k@���_˃���e�E�is�}�4T���EѾM��s�M����%������K��J9��mP�'o���Ч�#gƮ�ˤ���<"�j�B��O��'&=�<���	S�U� �C�)Rt�SO�����l��!�;X�(w� �n�68�7���9BW4c<�T�����,��h?��=�g������`V��Fɺ�ƯB�Xc�7XNj�4 ��{�kڤk�1։u媿 �6$Կ�"'t��a\E/��R��lԛM �W�t߷���p�ÓY/�����,��&N��L�3��vX����0cD�VE^s9�qk�Pl����4�E�9d��cğ�#ӥR�L���-��դ��$�T�����'V#�
a�ޯ��������v�t_� �B�b��_���=�e���įA�(�rLU�M�D�2����׼�ʻ�F�u��i�� \"M1�4�$Fe�I?����@C�sʰa����+���:��V3�K2j�ψX�H�`2mۓu�)��I���R<���ѕF �,`���ayY����
�������.��Fh"��NO��y� @��m�i�
1����W�&>�@������*Mv_��-�JSf��)�ᧃ����������fL)'�9�z�}�[^�7q��� �vKV+�Խ���Ө�E��,nt>6��0;���tj���}$%��h����g�X
[�`C�#�fd��;��E�"��A��)��HZ�̴?��w���-���A[��Q��,�ad�rY\-�����e:g�p�[��$ns�i����Ʈw��[>��4`CQ@\��g�x�-��4<�5��\��N��L2]��L 2��[A ��[1_��۪5��� k�@)�C>��k�dW	ԟ�3�e��{N��a�??��V�����D^9���3���F
+�W��I�7�L^\G���O�n$1�ٱ�Zu:"� �!�����$��#����� �b�&T��v#0^���4������'C�&���ۀ��e��Dq�:��;ǭ���@vU�֯|�U �7�X�bZ��%��4R�ӯ���_�N��#�w$���D�����q *d���a�:DO�q�B<׳r"*=a�":�!�.���}3"�9D��$h�g憓m�l���S��h�6���Fh��C&N4@�����L�Ô@pw5?#d�"���f�2�* ᫍ%�R�ӥ�Lm�����8LO<���2��˩d8
���E���	׳�h��φ��K��IBד9��� 0�U��m�Ţ9I�12�!JI���]dH'�""5x�������1*��M��sjL�_+����������Y�Z�,dj�x�C��g�b=�����~�u�����4�_��R�2 ��%Da���8�K�3s����ߴ�\?ڇ����������&/��и�;�_eP�w�jY0�d���{�
�~7�ʴ��콽e��R���4w���{����(ơ��*�S�x����y� �I7V��4Ev��"j$�"��ж��)�p,�i�:����I^�N]���!1��#��L�yj�|�(��ne(�A6ڠ��y� ^���d�����L�L}�q�;�U��Q:�ӯ���G-^��u޷�E%��
��w[�Y�0DD¯�t\?�4�>��x{��=T����x)�ۊ����GG�[l��������ta����A���n5�2|���<r��i�S9[/(��k��^s^y\d]���$��0f�hO�ʨ(����@���]	1���r}�έ�l9PvĐ�&�V��
�w}ş
u����#w���loG�#M�p��z��<HY���ᡗ�V&�ޭU��x����*O>w�v���>�Y���Ю�[|F���_\�N�9P´��͝�	�c�/Q�\y��q[>������դV�(����*+稻�7U��*�$gA��M���[�uݧ��s�E�,���9d��͌�W���'Ìc�LH �J5_�%R�ӻ& �^���4Ǧ�w)�ם��qh�t�s��OBY]��	��lr|������{��wiS����VM>�=f?N";�ɷAe��]ptd����|�K���/�B-0��uЈA�6`���4l%U����&#*�W7\����j�}���0�k�*����:7��֮͌g��OU��� )�l\[��Q����@�3��F��$�{;��G��;<Ig4��j�b
���R}�w� X�RVʚ�/�ՒR�w��&l�ƑK��#=�o��"{��p`=�+�������E�]7��<F�#�Xd1�Ky��1F$9��O!9��%_H�Y���$��{6��J^�x#�h����g};���O�/8��n�Ž���0��"�1�8G]��A�{5���?��EVm�H�i�7��M9��X.����``"��7�m͛����}��w�]u�������_�	B�ʱ�Z+���̾�䄊�<�0��i �T���{�5t��>(bC�JD�]��I��e
hC��8r>�Bc���
��T�.&MYX�	��`�\�|$=���ȗ���� �T�Q~!4ŔҔ� �ш�Ӳf�-Ӱ�nH�� B�_��v���^�欱-��B)a'����:���D�_Ui�gf>1qj�G�@��>~K���5x{`?�iR(T!�q�*�+b������SD1���L���'*�K)��[j��o���8�����R$ 5)�i�L���q�9^�ݡv|`����6f�օ�5�9Op�r�0��E�ߔK�����~K��<�XA
�eJF���˷EʵM<3D|0/uq��z�����dTJw��� ��D��rW��^���$�,~��p�a(���y��ԏ�T���v3�O���E�iB�A�H�&^5Y�Bn{���]�^3�F�V��?'���(~.OH<�/���1�|zn裰����ɟ^ܹ�U��"5�gpg�K_RL� @2�欩 8����cR���C��&eߦ�$Vr	ppB������"_ �pz���@���S,���l��U]X��5a�y����3�_��9���=�0��%�̙�K1z:j�nL"y�"nG�/1Ӥ�� ��\�=/@�����jk
�Y}6�
����;��ܮU��
�[�H�w���
���y�z�����p<K �U��' ��
�:��F�3��H�� �Ԟ,:����8���0�eC�@��L9n˓�◂����7��A�:��ߧ��!�Hx�֙A+:�c���s�?��7ʹ����oX;��L�1�f�Czھ�Ǔ0sf2�G�<�Ś]m����#�>����밴�}�S!s:�r>���^�ƈ���%�.X@��%50)�J�{�:��}lsa�x9cu�~g�f6H��1���!
�Zm$�S�=vo�D�Rd4�<�Z��)��P�a� �^�to���yY&ﾰ ����XgC����=��ڍ�XM�,~�h�>�:�^u�T�7v���mx|�Y�@6�vʳ�	7l�x�a��>U��D�Hȷ��}����4�xiO�G(aC��91f�+���|�y�a�lΨ���+z�1���.D���v�b����r@��G^ҳ]��Ox���}!��$7i<�:�h&��G@���S�ո����ǯ��o;~?@�>m��{)?[�:`}�����/�����69NCk2^T�»����Q��F/��ϹK^���������Ӿ�I[i�\0vqY�V��A?���1>�rR)=hk�~�۸�0�����6�z��<c�~	�~u:�|Q��)£�=c;;8�v��Z>�J\`8���2-��m����˫[�g��>(��=؍aZ���!d��w
żW��!�^E��E�WI��_�e,�1$c{�R�dR�MNOJ�2B��-���3�<��X�1/�gi��8ԡjt�-�;��uP��J�^w����ec��	�Hi[�������$�G���(&^d�]��E���>Z+H����˶x��Y'��z3[S�	(>���sC�}��T�UBx� 혢�;��x���gj���%�� �.��B5=ex�h����*?v*��˨YoS�c?z��"K�����S_kֈ?�r�������BEt��t���i��{��	&��q��D<Ҟg���g\����3.�@B���l��r��ݪG2!�&�<���٣XPB8�l.�o�E �G?���ҍ�y�@7 ��l|�)'`���l��9c
�7*p�+r{A�z�A�W*J�RX4�4fΪ�N��w��Ѯq�� ǨL[���m,Ӯ}O�	��P^-�����Lr-ڜЈ	N!�5ڵ�X�\&t�k8*�G!��v��G�����a���T�& ȣ�䠥��NE�҇˞kLe���~)[�\�o�*��,V����[��S��#�2@�X�@!h0�M��-���g��мi�7���-/}��)BKT�����`�9�x3��pǧ{~Q���Lh:��s_[����)K���!����)�4�0��T��z-���!��� Ŀ�������@7E��8�G`����Qly�<-�'�[�}�9�'���VQ�UQ�\$e���kz�*��}�W��0��،`$���h��_��2��'�����`n�KΉ�3���X[�_��@���~��Tr����=}���l�0�M��}Oj�=�;u��$����YA7Y�\����r�z	�8���l���d/�����j���t��<�_М�:���^p�ǅ|�a���ПE�8��;�Eؾ���A7n�]�|2؞���9���jV�r	���6#��3���;0��~@�E�B�&.d��(�N���f����q�ǽ����T��3��N���./�|�^ȸ�u���~�(߃�4�ώ/�� ]�� �ZI�48�pt�(C�*P%��?��i��P��� ���fe�>B�M0�=���f`�	%�!W!���􁴉�,$"�p&L1.�M)?�N2��uN�)����EMcl��+����}�%��,�;,��j�n��@V��졂� �m��bC��|G�nYSEװ�\vS%�H��MgҬwd}$�W �rҰ�p��H���{1���C�\��tO������`GA7��v�W���\y�c���?�u��mK�
q �����L�'{�V֔W8L@��^�-Ŕ �Ȫ�6Dj)�s����ծ�o���s����܇��FF�09B#�u�I�^�ݩ,69CU�.)����iPQ{?�u]�t���C��(%�5͹�R�:�}�i�5Q��>H�up�Xܢ���jｍ��s�6�A�5�.� &�!���C��r�n���{܏M�՛�5"Q|�<#y���XG�z|2��̀��)O&���'��PC�F���k��R(�A���y/�!��4sz��8�w��TU~M���,�#^n�8~���'���z������&��e�.R���K�G��O�<��+�~��4�����;Z��l�\*���d�D��G�B�|s �gqG�sc��C�L'��� ��7�E+v<�x�ǜ˾SћW7F��|�_� ?���l��8xd&�l���LgߛfV�nEg�S��l&f�ill�lre��]��rvc�M�J�ɻ�)���m�mFy�� ���Q��h^��Wv������-������G�r�������O��H��ᔤ�=�>k|>���ś�G�Ȍ����.$����pB�K�_�Ф��H�]\�)C�yoG����B!�����	�H0<;4����7[����ZD��_� �-atH!������)��#�W��+mV�CD�&�P��)5��@�\_���]�QO�� Ja��S��73����d��\�}xb�؟����\LR�8b5��+�$�����QI2s�`%�,��K( @�c�@�_y��'���rN86�/�̽v��|vkvh���X�#|^����H��Pu�F�}��Z0w��KDip�ۊ�^�QE�'�'H�ca��
cg�T�kLM��$���e����/�Y9g�~��RR:��<��d�������^ +���T�q2�L��Ӹ����`��}��q�����2[.��v��tΨ.�c���ߌ��wM�z�T��/Sף�L���a�5�0
�J�I�%���J,��#��'���+(�.ƀ���D���Ol8��<�&C�d,���>(.�t?u��ݦs��2mm*��OG猶\9S��]0���a��KxM�[_��?݆�$�(�;��*�T���������3�G��V�����y���"ęQ��F��~����A��P�0j�P� eվ���85 �H�T60��oY��-�����
�qY}���'u�A�l�?Y�Ái��#j�H<�J�SH���-�O �\dO�r�z�}��P"5��i�ǰ���Tڱp<������51��_=P֎��e4&��h�����e�X�ߘn+A���wUI�5;isx�f�@���((��0
8�ˇ���ѳT�