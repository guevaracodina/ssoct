��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ��p"���C��T�fX��k�+��)��6�'�3��$���)��2�+�
�#�7��Ib����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^0�"������֦g��'�Vv����qI��C�M`����⢃��c�
��rH�pɡϊ��0^k�?_	�̢%�1�0�ְ�>I]�;�걵�s�i!!G	͛�k;gS�?'���(�|=a��!a�dRPP�_��ݴP���C���u�)\S|���_TB�5�1�%���̽In�-�oDx��>�6")�KQ���D�Q��n3.���n�)M�:�h='h<���:LuM��[�A9�۷Yt<Q�x,",��9���^Q����Y9���n#�!��$;��1\�9�!u+C<?�P�_�U���O�Wm�+�!T��VȎq�tR@'�7�3!y�С�@dߘT�0AFEaIY��V�Ǎ#�	 X�8Y'�gB��� U!����xe�2��`Tc��^��>�Q]���֣wA>j�+�: ��9�b�!�8 f���+.hפ��}x4w-�lc(d�Ya~qu�k4 ��CK�˸��t��F���)�����C�Q���X��Sc�
�������?���"�c���[�N�[��b����mqB��aסA�X���r(TW���}�U�a{��g�O ��DD�x1�˜��6��i^�ʋ���	�;M�L�Ǘn�����R�	� $ ���x��� d'��1�F�C�u�w�&���W��Ǔ�[E�qk3�7���n�>I��^��.��0 	�[ᓧ���/Yz���o�3�Q�Rn��\��!����^��ʌS�P׃�(o��I/گ�w.ǡ7��pI�SC�P�=����Tv���d"+��jS'��Q�
"����Y-�������&�uM�_��3W{i�(ݏ�����`�k�d�u���ո\�o"�w����X*�1�Vp��C2�:��L��z����o�A6�%�[ӵOe@�R`�+��yZ����z�0�:��gɮ�����Q.��\�j������X����_��<8l԰���=�|+��&����[�k��F7,�7���^䴽e�t��$�?��8�?Ҝq�L�l�|{=5>{v�K�l���G:��{؃����Nh�� 69����d�J�~XN��aڢ	���!��W����2<�õ��W2�_�~�'m~	y3���@r#m�-����n�h��g����/��˸����n��%6H��MY�.ś&�s(Jw$��@hr��s�����X}��$�Q �-0�r���P(w'�8 �s��V��ǰ���d/8&V��!�����Us�t���������Re�#~-	0ԑv y��_P&� �a���}AϤ(D:�.If��< �������ԊN۳g�9��9ΰy�SF��^���=2�`�,��t��f�f��4��֠:�����p��T~��l�Vר�W����Mr�����j�'̉L��^�;��7����	b
r�ߚ��`�y�'�(A=*s�>�#1C���r��ʣ|�:��&e?+�F����yWZǄz�����1�[�>�Q	������R{�TسM�f
�=�_܁1��J(�9Ns�YV�/ ��3G�M!�x�'�V�f�K�*f���]��B���J0��� ��}Q��=��gE4���cR�M���'u��t�j���=����3+?�IH[��V$�o3+sWϽD$��q9I%�8��O�S������ ��"}�ʘm���Y(�YKG��ؠ�����0�p�`��0o�X�_
��'�|��U��l5���i�[�6���iF�W���^2։�|SsgdPz�8�N���~�����3Ƶ��f*��;bֱ��\�����G"��;]R?�W�k�j�3+�]<��50���X�4Jlix>�S*S�T�	N!��<��8s�4�Z!�[X�>{����ᄏ����Eo2G،mҧ^�i f�/L����-ĺ-������<�s�qskx���P0���c�B#ơ�>@1�'��BG*|��G�r���!�Gf\��j�_��QE�%��c�)�rESi$nճ;�'-9�Ne@���<P�'�N�0�d�G�.�n�[kF��m�'����(��||J��%�1=2�� ��5Xf���B��T��?w�PY��k�z�ؐc����_p��#e�E6��U�a��C�	x�o�×!�^Ȅ�� �O	����fN�^V����`MɝϹ"\��ZB�2cu9*6�^t�*���L.0*�Ɯ���ī�˷r!��� )��:GHL�`�7꧿�ON~(��8r�����ޝ	H���@1�e;E��7;�Z��%搅�	�:nr���?�\̭��T8 �^�6R�֬��8�MYgW}�vICV>=򩊫j�dk�f�`sP5��g�iu"�M�\�:a��K�U/%mn ��%�5ɥ<��,ʴ�������L�2���;�%�~x�[��Q�8��Gr)Keg���,�W���-�ɪ���?M/E�ph��s}v(�W4"��?I�2HȻ;YS��{�y���.��]�YX�-�W��D�"�~c�0 ����g�wK�KC��z��d�� �"G���~@l��X�2��Ȏ� a��(�nf��k�����K0"�d`r{����{���,=@� �.2	>�Ny|ҮܚAue�^n I~�ٙ�ը�3x`�]3%|�P��6�[��� ��֧K����q@��$?�h.PW���d��_�S�ZU@�B� @�޴�',
��⇓�5�
U����e'B���)>��2�%�� �92�7���ԟ�U���cХ]l94y�J���Rj�������/G
"��q�۰eY���4���H����Sή��m���2�2i������W@���MG�Қ��ܷ�9y7+������ս�+��t����:���R���)f�����d�c��Y�Y[k�sb5'�I�M�=ڵO�����]�H�$Ȑ���~�@7[v������S~'���,�e��Q��'���M�l�ʆ����u﫮sY�N�p+'��6Z�7z��9��
t����*6R��ű�V�t�N�چj�n���AFBY���@6�}�����h����d0 �
_��*R J��ڥB�YJ�,�qlL���U��r��O3"	v�e�m���P�򵏝1��j���ie@�y{t�b0Nx)�Y�U�P�.v�������}����}>����'�B|�{ZvaHw��q���O6���~j�$ ЛA���� �xO�@^��'�j��Ҽ��Hp����s{���
u�\!�F�e���{�4���=��}MKc[^�`��jԃ{�\���դ�˦ �(a�'����W���.+4���P#O-ט����ɟ���fd�P�cu�6g��XQ���"Fэ6�!g�l��A���yZ�+� �Q1��:�^O��4=��1�mGAn;�_#4�v��p�����h'��c��H�����ڹ��d�a��Uw�؂�*�����0��5��+СD⳸�~8�ǢA�q�$��|JP�o��K�=�5�m�Q�(/N"\C&D��
� ��[��t�+M��}�����ay�
PZ�	��_�bJ�vl�Z?q�sW�#�٤3-9CM�=��)��L}��;^q��1�Uk��,C�Z������Ӈ���\�����8�8q.�%Bj� t1�N�2��iw�py�4M��c�G�#Iw�@C�r.�J���z :��hv(]h�8:��kv���� ���)�K�~TL�֯Zz�N#Ҵ�0��,�=L�Z����!Wߤ�>����S���^V!��n�u A��4O~�����wq�jZ`p���s�͐N��ްW=8� ��V���?o=��<��e](��1�	[l��:t���%�8J�M��
���4܋�o'�!�yӤ�c5SIY�.L�_V�1ͱ�g��ޏ��3��-9k��O?f�y׉6�����%�^l{��{�?�(I�"&�vp��3�M�P�߼~束|�w�'�Q]k3z�4!�x�����w��n��S���WP���g�֊�� �7��\��z,5�F������<q���"_��碼�U�lr�,I?����)� �CXz"��ixv)�i?f�W�m�>4�=��o���9�)�у���5sc3�2�<3�<)w��&��H(���\���P�݇NR������?N��|$�y��&�'����B��~���^���He����5|�t'.�	'�DZJ�Q�ёq���! j�G-eNcNe���C�c���1�%�5����(�je����?�[vDi�2�'L�l�EL�o�?�w�l��6�m�ɌcCz��[}�c���<�,N���,�g�Wg�m���K\��1 �rhq�1]�q�{K���X�����b?�FK��F�]"I�4��s.��ː�-���[�و�ftl?��$��^�@r���Sm\K����9�=�uLʆMK��T,۠󑺊S66�L�s�1�_�����#8B�x�{�F�{R�2��<2�C��������J�0��'`���Yx1Ky�B��	�q��g�/�b��1�hdQŒ��_^����U��'���Bٓz��.<,�2��]��#T���S)��e�L�H�e��(R �F�v0B�����2Z�#���#���7Y_(�h�K��QK%vj+������M|��j�O]c�0��IT��y��4 �ȗa�L9� kz��g4�����:	���"��XE��C��.��%�.����Z�<u�P�ZlU��s����F�$N��v�	�D<󥩕��.���6�T��λ�d�n��t#k�Z#���XQN5�Dcm��`��(B%���d��þeu(
gC�,�!�����j	|@�Ȭ�x���g���<���#��P�|�f:�՘��'؍����ʐ~����sw��.������vm1���3X{�1�C��i�AqX��՚I��y��R]ʎ$��h������z�F9���]J�P?+�g0<b�oNƺt��]ΪJ���αI�X��$
غ�f�{vX���X�>H�ޮD\ب�	��?��� �-��%l�C�=�d�D�!���f�C�=�g.�_�y�i��:���b#]���K�5P�!��n<E<�T�S�u-U�����cTH�\���q���PN��e����լ�G��>�M�G�g^xr�UQBHr�u��ۢi�U�ķ�=.�J�)�Sa����	�;`i��8�����)�^(v���FC�s�q9gRuLX-�,�r��Hﵪ."��k�k�@�I&�Zꮬ���@�jӏ!�
@�,��yn�@"X��W���9�Aָ�Od8���p��x���ɾ�$�ʀ��cX�迄�#�qc��JEj�X�.R	�~8 ��k!)*Q�#\z��]d�c��9�T�/N�iya+ݷR�N���r;l�x�q��%ܳޮۉI
�]"Z)=�g��xT��ݗ�/����Z�D�J@إ�ٍ�\�6�X�"=��C�J3�`�@��㖕��(��+N(<�V���l�i`��4q��P=��&��~͹�۔����-drU��P)�l���QQP6�vt	_a�W2�Z��:�Z6z;{�='y,o�r4��FyP�I�'�|�F�O ���J0�%���8�«�p��[X���㞎�D�ƕ>����kL�
����k|��[Z��]�ݕ��˿��f�@���y�*q�Xy���9<�)���2*ٛ��*�۬G_�#�Li�*���r�݈�K����9�����u�s�;��\bn�6l�BV��ˣ����z| Jn�KGȼq� 
����\�'��0x�e[ O�v=�da���P�S�x�8�O�y, _e����߀�9N�ū�!$M�&06��f���>��_]�eHc(��D�����I��\�5��Щ��Ē���,�f��A�i�Q��}��<�}�r,��@mV�>y�\���2�����|�������Mf{�-Bź�҇������؟��L�Z!}g08�=x�8�u�+��3x6����Ǽ�٤���tI-F�?�P�yGDב�ϵ ˃�Mg����+����5T����-�Ľ�!�)E�{�
����$�VC���`&{�O3|�<·Hx�/�յ�a�Q�,�)����'_J~���U�.�e�ho��{n���i������ �@Ȫ�v��.�ܭ7+�a��o�Ϊcy?0^ �YW-Tdy�8�GF�h6��	�I��w*O����B�U���N �sJ��Wz:6��E'M������b5t��@F��V�p"�:��vެ/�����GGu'� �	������%�_�:�\��u6A�gJ+%4w���T�E'Bۯ}gvQ�8��o@]�;�=�H�o��.PHtާl+�%��!qn��)���o�tcGw�	�.�h^n�1o�< i-��egE2��c#����8S�[nʐ�T�gCي���	s�
]o�aq��24��3����+�z�&��a��$TM�a�[�
�`{����ܖ����.��7�N�^�,���{b|�P!�)�� �i�=�d/j�=V~
g~귓�͠�5��G��L[���.��g5Pt#�ܤIѧ�,�	-��Ϩ̈��S/һ�3���E�ȴ��R+�6�y�f>Q_m�&�b�oq݅���t��l�(�����c�����[p:*��n�E��;0����2������n�W��Pe����#�_WxYjL����
���;3�L	�D�W͍d!�_+h���9�[O��$n���� ??z�:�И?����y� x2��Z/�wi�}�~�K���@���q��^Ê��V�s�K.�3"����o�9i����2];��<���D?�H��������{+���*�|�l;���5�wp�	�� G����s�e�o�tx&)U�cw|�AoX+���񊙏�1X~��� 	�Y�ʉ��t��%��Z^qJ�c��",�y��_��a���<�L�R߶�__c��y�=��1{uEG��7���C�b��d�ذ��k�����T���?�g�ݫ`�	�I�C�!n��� ����9�2E�)8AĽ�nN���R\��<!�E��$��]d%#������<��D;)�:T�4QIJN�����ͼ��U&����+'e͐�إ/�p�W�h����_�Kϥ�H@p�EOOT?A��e�D�QKnw��Z��~�⇁yx8Dl�C���+����4�9�Qd����)���\���}/.\���D����H[˩�s��ǻgYQ+<�v���)�kK�Ik7��)8���2nڧ�7R�
�� cJ��wպ��E��YSA0zZ&�-�G�K���-ȿl�b�$(w5�sf|�Q]��gc�u��ʧ}i�G^�݄z	"	7yB%�V�N��{+��YC�����R.{&S��_��=�����V��@gJ0����N�EY1[�pD�����.ߺ�؀���RX�C�X��GG^�w:�f�LGpR��Ŝ���h����ͥ�ʄS��1����k�LZ��/��.���՗��V�2��[>9��F�
a� D`/�y*b�ⱊk��%�(�O/v������U�F�O�*������a�����X#ӱ:5{��:/�؆�	�u�GmdH����-���f�{N���2nN4���I���ni5[ukkY� �y�{u2�lj��`i�tz�N,��}�Q�+�T�_�
~*)��j��x��<)�3���z4`���7��;K�!hur64�����(��Ii��2�D�>�G�c����pB+ho���H|9�DĲz��HۉJt�gQ$��^Pc����@�M��6���uªyaح��'YaX#���ӷ��Z\A���#�;*(RF���r��B�`&x����z���OT���d�����I���8]ѷ�b+I�ɬ	�_JJ������@`���6���p}#�����Y��~Y���"��U�0�z�I����7#EQ�0�?�9�c,�2q<b�rK=���|���aHAl]5��x/^�#TZ�"��%6{���~C�ɾ#��b]K� _�d�ǧr�?��2s�!���Y��4��^E��-�j�Α먨�������ig����[w���L�w*0����a���6��o��[]��~
����^�>Xӄ���ŉ�D[���S�����8r�J�.#&o��>D�U��@9���);�F���#a�A��D����O�a��k��z�׽�����fc������~�P��Vv=�:A�c����,��jW142�k���d��l�qm9����s��#p_��h	�u�d� ��<�}ɨ�Nd]N����,�!�2���{�lU��Lx�5�@&D�wAO�k�<�-z�)�'zSڮ��ͮ�&îHWB�ը'�$x�����v��<���|�Pq��!�=���c�;��THT�u1J��[�j],�+��9��G\�[<u��d}�F�Z;)J���X�Gdh����:�8���,�T��&[���-����n<[�g"]�����^�4.hF�V�ݧ��U1���ՙ_~̗rѕH���M�܏���^����P�k�	�o�K}zL\�o$R��m ���L"˒��@P�c��׍�Y6ɵ�*��}�	0�l�QE-�Y�ud� �d�C���1 Á��J.�,������"�}��\i�Jn�h��)�,Pn�Er<b�()a�<�[�A|����/���3I�dlh@N�5���w@�6z��⌬��3ؘc􋌳R��y1Xkl��W�H;�9�.3�[ �=l�a�RE�II����ۣq�[	��^�k��!^k!~+J&�/2Z�vb�u����
�pɭ�f��q���q�T󁬢�xi�c��lka���|#�� �p'���� C���y��`zU��գ��獵����W_6����Fo	���gt�D�l�I���[�@ē'�޺H�K���.����Ǭ��D�v��q�^�3��)F�;^f�B8�p`�v8LN��{SM�Jz����s�Z�%0ȡ�����gR�z��[�X1&�9���+__���}�4h�)�0U����l�RnFy���Pq�� �Q�k� F~�Tu6�&�%#9k�Ѯ����x�1�
UH�H���]��y���eԢ<?��{�~�g-B���g��B9߹�L�^��d_�>`����K�UJf+E��(�ɰ���4�P�)հ�L��m.�A�sP|R!~�eԍ�L{r�>x��
[���``�~[�&^
��m�@�xy��B� ��68`��'=欮b]�o�ˣ�؇��Im����Bq%�HF'�\�|W��S�tq���{��r�+േ~����@��a,�����2	cm	��K�>�>���5Xvn3��Z��w����&l悑 ��\T���>��0}���5�H_$�W�,Wܘ������~���G�ܝ^���� ..�W�����ƒxC����Y�(������μb��/z����ȇ���Ng�t����=w�sV��d����߻�Y�l�|�w(��.[�[�$n5~#ބ��`E<��'�n|���Po�+�'*mȾ���;�b�P��9��o����(gi���YJ��T��ʼ©�p@'��.H���j�mˣ ������+���˳��r�`awN�p��0��h(D@����CH�a�����,Q��x�8Q.@�/���%A�ţ8x�\C��h�
#��ܰ���x3��,��εOi�!�Q������4�����]��Vq#��}����l8�=x @�>	$����*������^��kBQn �xf��&QYQ�T�ɂ�<�,J�ݦUK~��y%�Dm�h��$�P���~���)���a
�y/�*�S�����uQ����s.���:\)N�y0]�W����� �|M���Nݔ�O��f�cc��Fl��.��I����]�"|5���i/��X/�h��u< q̫�&b�m}��e���a��Y{���`�	4��쩯�x���D3�b�o)eւ���k7]'FEѾ8�g���G�CB�8�s�Ƈ��=8I�\��8c+Efp?O����lf�q��r����"]=�s��4�ϥ`_�1vpsNgY�I�C��(��!V�Pυ��=���c|��������KX�3-:n���OR���2n�:����E�d�@o���t`��o*��i�������P�g�0��F�k�0�yF"��x��h@{�q9Hƞ�o�ތ��穬��n�o~���

SH����~g�֨� ��s��z����7Z�����D}�|&!���f�R��o�cr\�a'W��G	B��VH��o�]�Y>�}p;@��2���D�w�	p�'p7��ѝ��	P�l�|�_�4��)O���!>����\���*m��ZA����Jڠ�-�!:N�O3hȊrU8���hDМxG=����y��|���JW��'�iru�D��^����o+�^�&xҎ�*��W��1��3�,��eI��L}#g��oC�Ј��+|�dڒ�0��J�֫Z�b!	��.�h�N�_�h{jwR����g���Y�;< <T๳h'�L���C��>7	�V��Jo�KӺ"��R,ȫ:�|�%̶>m����ֈ�h��e�tB���N��dtq�cj<~ƶm�U�*%��g	pM�^irߺ�Q��Z*F�>q���ո+�5\�jm��A6/��n��0�
H;�'[�Ԓ�eϗ";f<��n�YD�ǯ:�l�xIo���/@�~���x�#{2[��v<��)��[��`@U2A���p;~�_ �q���\�tE�������3$QU���G�ZB+O��jG�Q�A�ά7�^�QB�iklGR1)�4�*C������ܵ��i��Z,+�wx����+��Z_ʜ�0g-n=����]p�/�(�/ED}�/����=e]MB�=����V��Y�L��qP�{ҏh�氺�9��tO'Q._�&�U �Y��?���ے���;�l���ՒP/g�x��H$�s{h#katY��P.c����5>��>AT��ƥ�Ά(B^f��,[��cG:C�,o�E�gO�3�v�h�ޜE�X�<7�6���~y��U�)�Rއ��I�O�[ �K������N�n�#�q�w�E&�#�=���<Y��O�ҥ��������4zܻ�c�X}� �|j��ģm!"�d�;��vn���w}zt��=���ļ�!��
n��uHMv�<�v����d�U���M����E��y��B��d��RB�h����Lʍ@ Q'��j��v�g�/�3	�AQ4�w��r�=�ٝ-���ଛ ^�K����Df��!�_���N�A�d��o�p���)�*w��8�η��W�3[�
�.yX��T
�i`��~��
��|��h��,�l�I�@��MB���$�G���@����=>]�p��y�:��e'�����,b-�?�OU�];?�~O$�ؘ�;hw��k��'����`~ًYS�d:�%�y3c��
�Ҧ*9�Q�Aُ�`'t�?��u����@��i-�(2=�l:�mO�Ӭw�V�	JZ1�Kb�b�]�5:%!��q9�����o(N�s��b� zb��e0�g˪|_�qv�_��8���fر�H~�����bW�Z�y�n_ �$�FH��~�i��S�eTk�7Li�u�{];����cA؇TAۗ��c�w��ӿ ���y64���)D��qW��]�}�n�-1��l� �L$�����-�>�A:5����#�7&W�##*A��v������0zXc[^P�\�a?M���#fVX�[�s_.`s]��uX(�ҁ�oN*�n�{`��؄������U�WM #W~À�a��mW>����:>͊�rS����~�8JT�ǎ��<ʓ�0����� /���˱	 )�&4�=�];h.�A�b�����lǵ���0 8B
�����"��boVQ�E�.Oj󅄚�j��,��/�b�i5�z��f&�g��@��b��S�O�N� хg<��W���P�'٠&�i�/Gt�o�F���돑��s� f��=�Xn�V��^�.���(K������ާ����=N��;�"릗����!q>���P��!|Xݍ~�6������+x �|��I��b�����F��������l�nL����W�G�����<6���6�|홽�(���~��ϐ����4��Q{�G;b�U��CK� ��
��|{��������D��H�.�tv�8W��~?�+$1�D���:�]oӰ@C���Y�u�� (P��
��ESʾ|-��{q�}�4%��$vB��gʨsi�r�5+X�u��%�����'n8B�ve��3�W���X�G�K��^��h[;7="������O b��'(��`98�M^m֋;��ɳI����Iɣ������!?q�g˷��`���ӛ�Z�S����*�"t���皦�M��Ukt��W�6!}��`�k��j�&:�Nr=�_��`̎����@�괐��\{s�H/��Jl�<���,/'U��A;�e�1O11�|����1�͝��Vx����;�(`���n�dJ�>����+���v��2��2m�ĵ�l�C_l����s��A�%���Q]�O����)�/Q(��A�[J�rvX� ���|��`��ۻ�4����6ELc2��-B�̼?��ѻ�1Mt׍{Ŀ�~�5�U���ӱϠ�?�&P*~��-�A�sN��bV�ׄ����ƏKJ�$��hjc_X�8,�3�>��$%�,t�UmԆQ ֭2-�55�O��\crz4<rF�x%��gT���o'!>�f1������K�kCD�~c��!����5Ъ\%�|��A��0���<�IQ-:ñ�d�~hH�4����K���6)�g��ϱ	}�Y���2o4/�����s�|�s��HE����=���_>��B\8��MuMS����`�N5�$��VՌB&B_go��{�2�c�c���ҕ���r;��;'q9��H������]z_3z_+q��ҳ�.�8�.��M���ϳa�Y��+G�+(�u�V$�|?�v R���B�Lډ9c~�bGq�z ������㴵�{x��軮g�?�Y�譞���2e�Z�$�o
�x1Θ�(�𗳟�8�� �:	� Ӽ�}\�������w�6��n���fW�P/�e@9�GP �
��9Lr �!�6�Nw7�ݬi�A+����G�ܙ�t����Y�Vѓ81��׳n��$�����8�'�P#t��9�`��^1l�1�	���t���6B�3A��չv �_��p�Y�7pԆ"�4r�<)�wh[��K8�7xV�� 8�w&w1�Ж�mFa���b�\�tԺ�z�zN�W�[�F�@�q;��nd���
f���A�#�Y3���b�a6�񭤎e���F�C����]�2ʽ�=,���|�����S��<���	{K�Y4R���/�%b��੧Y�Q��2X�4���G���ʘ��`K�\��_�vߘ:��Jcjśi�ʔBol(��wgE��'M'��^`�W�^����5�:9�?FS��5j#Tw��=V����kI!`�����PC��wǉ��
&^�A�ZK��̙]�Q���)�J���_��%\15\��讍�C�/5�.����|��K~,v�2�cz7c�e�&�I����
���[�N����sz��Vqy\�v����'��R���j���j:������2�KHɓ!�8f�P��]��$�,8K�q�^�/���iU'�%i����J�g��!}\$�����h�gf����%�%��z��Z��ΖEFU.]��7 rL�t����AG=�;�"��9=���|� �ʾ�D
I�O"��:�S
S`Ƥ��G��ҝg��'#�T^`�����S��K�W��΍^�wSZ�a5��ÿ&�ڃƲ[�h�R;&�����0Ĺ��ZC��� �Ɇ��o=��8O����e�؀N�LSO�@���9Lw�����X��0vnE���GrǥNA�?�b+��p9�5}��0��sj�}�� ��:@cI~m� T�;@���:I��)?��X5|���.I�6El�[��KX��� ��3~��8���ѶR��A&�{��/m�
p��կ1��t.��V���N�EQ�,���9]������E$!K���E�W:�%�Ԓ�cmO�F��t�W��G��,Ƨp0[&�?ħ��c_�,6Ho���Ixf����+�U���_w!�a�g��l_rr�� *���?���V���\�b���\���r\[���R�$�ǘ�ߔ�\�� B��zlL�Y�K��ɨ4�q��>��g\�a4w|˘��_Ɔ��O�b��S��d檖@����Z?��c^l���]����e��q�E�=���o@�
���ѐPo�倖�h��ՔǪ�g�� �ڑMJ<-ʅ�+$'�#vi���X�~�����48`����!I'Ġ�*���:0�8g��瞂����5|�9(SG0��'2�|�����?̓����[��%'�A�����T��N��dۓ�uO�����:�Cw�2���3�H�
�Y4�r�̅5&c&������ٸ��񮭂���#b|Lv����7��ԲI7:��Ff��<�]�	��*K���Ѓ���gY5jh|��-�����œ�$0��=�{��5��e|�v*ʣP� ���%�9ִt�nǖ���/R*�U�ҵ��o�l ������s:}���)��u@�1����Yl��BF��0cJb�����v�&�������եQ�1�#���~۰^������9�h�P��ܙ��Jhg�@�E�O��tSt��Abh'�o�=v&`�!���f�#G��,��"�k`Y�\?w�S*e�t$<�߇������9	�v�^j�pD�"~�J,O��i�{f+ P�7u-!�tA-�8�/?D�'U�o>�~n,u�>�����-�;G�%�%��%��p��X#���dL'T�,��9;�̈�rȸ��uw�>Ϥ�+X�+hi�r+�/>oo���Em�YKV8�Q��XI�Ą=��r���C+*Mw̙̡���t�|1�6da��_?�vP�QB���a�Z\�?,������:�����؏ޝ�pF���^���p�}�e�&�%�����e��QbX}�M	��F��H<SP��d����]�	W��?�|�Z��,QM�M�*�#Л�ڦ� ˑ!G@�U�1�����M{�`g�9ɴ�k��JG��湛_�q�Ry�k��\}|�b�Û}�y��YF���N�.[�K�)�u��O��#-ЖzuN�,;l}��>�B0����+�u�ٱ�°a����� ��Q���s�0��7-p�R��k3����Z��P���	�t�$*�F}먻�=c[<��S˖���0��y����f;6R=���,�+����{q�숈�.�\����_�t�b��f�5AQ+��m�\C�6⾋�J�� ZV�K�a�ɩ�j9���� ��*gZm�S�5+��d.��{�^�5�c1��j)Q���hi�����d�ޅ��qۊ};{"C��s��)	��4�h�x�m"yH���$�=Xu���c"
fp��� �=�O�V�th>˛ب��~*hȊo��ǭ�]��PѶTY�#;˖Wؘ�(�	��2`gY��(sd	U�/�ɼ9x��JA����ilG���=�l۟����0�A�� �D��e�ɜY�i�k�@�g���\<O���\<#:��	)/�L�4�����c$�Ur���%�E�C�G��/�]^��=��U�"��A��cD�p�6H�iF��oީ�N��k.�M��R��M��t�]U����;ܐ�ba��00�����p�d�6hl�U<����;SB�x2�7pvDD�`�@ܺ���5����D'�f��yt�#��y3���0eA�4c���ܾf7�!ã0>�l��wjARDib�W�ŗ�aG@HH����!���$�dg�񀼆�vc��I&��d��%/Y}�N޲�;9��0�F���Z2<�.�=�*�ʡ����F�K��Ǉ��,�#���Y>]]��@SO$���an�סb�L1mm(��z^<�U�i�E�+*@^m7R�{�
��+�0�p�~+] B�G�"��
5q�`��c������ѽ]�b+��迏m�T�-���+��;�8��6a�j�L���� β�I�S�w��
�hs�	�}����������cO��d�t�w[���)�icO�7�>���S/
�-�T�u��
d���l;��f�ckA�ϊ_�6�
��1+���T������Ti4�8?%/�}H�ԴU�aN�z�J��Wx�nr�ۢ����h"�$�YjL�m�����TT���/(Jo�������B��� ž�1p3d���R~D��k�#Y�T�Q�7
k�O͔�n�������*^P� ���[[���o;�Dق�NV[�f9t�e��T�mkSŝ�Y���O���/��M��Xax��C#�n77�6\��;?��-���O�?�.OmLSh���Ϗ�-3@�׿W��?�����D���Y�5sYk�L�,��-zV�����q�����;2��Zy?�g��U�jl
��㔨�a��h�n�ϫ̡M<��=����NU��;߈�^��@�jL�zOE�p�W�!��}�Qz�mnGr0� h��N����[S��.��<~���n䚶��tsŕ��� q��%CJ�M���@\I�p�G��k��y����u�*��\
BeQ�\�f���Y~	35}[��ӱ�>e�L:��#�c���hn��oa	��h��T|9��D����/^��T��E��J�A������;x���:<�E�٪����Ows��q�d�+,;��+?`"]�\���i���ôU(Kh�ZIQ��w�iʒV`Ͳh�'�*�!���z*0�U��B��x��_�qB-9T(��	�ʯ��&��]�̋�ˉe(X3Ep��~`�_:A~��ҋ����Y���,�:C� 3wS��%4�`�1/d�����}�·��S���:��\�@�(WC�_O��V�y3N�oH�o�ƿ�a�C���Y���5�J�|��D\�	H�͍��_�����}*
�bp�qA�������h,�^2d�Y~�z�{EDR���|������fQ�%�dH�����`P�zf�y�m� R�F�
��)�?�y�c
�6|5�+v|pmwߞ��8C�[�o�s��x�'�G�4�X�v���?{��A0���
k�.��R^�6��b�2n��)uำ+�b
C�k�HG6>�`U��ӯ�Q'0�C�m���ź����c�ܜ۲�"G>�H�ӑ�ߓ�a�R��*�c�e� �t���~�rh��G��;���m���z�E�e�`��K ���ڻ޶-'V�ͩ�o����Wz�%*�U�46�s�0�{u��DbI�@���*O�mnr/A�ê*R05^��v���_�'l�2�`	�Hoa���?Ꮮmy�aW
�iD�NAI0�qc�^��B{���nK�H5��D)�T�V�^:gS�'�d���t��I���r���d6�W��ؓ�8�ُQ#lG;��{��o�pܺI �4��f�7v��V�nG��)�%�&�6z/i�G��0 3����c��%�O�Q��`�������
���$G6_�2��C��~�\�9|�	@t�W-��"l�=ue&�J�8; �	���d�AP
��PG� 3R"U�o�����n�O=���V@ce�J��+��ig'x|���3��\�6!���Q×�]��p�Ր�[��F�sRO(��u�����	��*+`a&�R�H �����/ ���A�]�Z����寫�E�H�h*��>P��d͜~���cbZ��nx%�ey�+��"\�e�d��zR����W���0��݄{ׁr+�3��,�ҳ5Rn�� ��{�[e�/#��P�:��`�&܉���ۏ��C��V�b�������M��>��r>��.����#'�}���-˥|�E�R���	��n�eq�H�ۜ�ھ��x��a����%#ܬ.������T��O����hU�q+�5~Z.[6��<j�"�#�(F���p��-�ne4������t�ǳ���?ƕ˅	�E�w��\�{� ���l�1��G�.���3�v/9a3O�fP���|�݊�P��6���ֿiQYjUJ���&�t��D؄ ���ڞ��B[ͦ���!J�W]TV��H�L�2ujQ��sT����(˘�`��ѓ��[�na�	��S\����j�y��5������,����>un�Y^h����d�|��o_?+�DÈf7B��z���G,W���]�\��w_��MՁ�3�qt7�5�3�\�bp�ׅ����d<�*d �ahUv�iW�^'WA��(`)�~����xH�d�p����7M�� g紱�7��qBg�E,3�7�3�{1@�o�e���Lv�$0+���{��e��tVlc��%ϝ���4,�2�0��Q�*g��J~m��ޑ6�xtR\:���o�M��\�j���T��+�6�>Y��rtR;q�:����C�FPC�
��=�øĳ��@(ׂq�F�n�Nj��0s�K6p�-�$*�����{!z�6~X�4m������3i�n{�x�W�� ���4�a�/��~9�?~��\������{����&iUE��	W0��7�k�vm��@@����P#��I�vH�%�QMJ3���J���*��ً�3��a gd�^g��sp�;��9�<r	a����"�-���e}2��Oa+B�6!�S�xK�j�uV :�S��j�˵"�ϨA��cz��_���� �����w�v�K���,�y]
AŪ"<�.��k���8jE��َ!���M�|�<tk"�U&�Q�|�8q1�K�-ƓN�$��H	h�����^8SH���j�2���S���1ZB�=K����XS!�=�ΰ��LV�1���e<�U�
��]ې,+��܉��J��Z&}~?�b*��6ٳ�Ă�̓@���dIa��P�{�8n�$�ۘU��SH��1�y���N#Wy7�̛��ט6�׿�F��K�)M�$MF��K���:�!�Y�w�8�G4~��^�F�@ez'�� ����`������}r�DG>��R޴`��Qյ�kT��M(������]�P��I�(�/����t>
�-PF
� ��!��Β�����g�BkzV�O\��;@?��{���������1�w�ר�G�ɹ*�gv�MP��vH�mQ&�4qE�lG��M�o��aGIS���t�~����
S�R���� ](��1Z.`Ar���/'�xУS�L�����g��$�t������^'����Ӎv��X�NH~?]�Z�����Ҩ��zw�F�3m��j�Z%�R'0�H�����d0���z�3O��7��������*���e�#��ޙ情�zI���>������H��偉V*dm�,�EA�C	0olRf���c�7X�J�	��1�`���
|!H8֜['}�G'ݫ��,��/V��65�ZY�	y� ��� *��~�-մǤ3����|^Usb�)8�Ͼv���Ei˝����_��� ����5R��\8p��<ε���}$�E�:T�~'�hoȂ���lK `=<������E�3�#��엤�:�l5i�\lZ,]�x�|PJN}�S�m�oS�{�B0��ԏ����j�����/1�3�4�^`�^��H�+���ؙEp�hRA:XZ2Scr�xz t���]ז`�߽rg�� ��"k/�R���C�z�A� g���2�s�V/�9��g�����٢��0KL�9(��:���L��{�V��F1z%����I��7x͟�K1i�,���֝�0<���]�М��:)�)��0��4zי�Jx�g(�`�qr��;x��:��cG�H�86���q�V妅�r�`