��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���9M�;y�f4��]��:��&���&����*۶?�H�ƃ��p"���C��T�fX��k�+��)��6�'�3��$���)��2�+�
�#�7��Ib����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ��l�� ��f�C�9��u�Xv� >P��Ɛ�)u���8�5�N��
{��I������k��RV �z��ˋ���!U��^zZ(�V����S~R4�~Ϸ�2�˞<?�_4o��o���
�
$��~H�BnѤ�Ω��2����:H\��+ֳ�Ü��[��bۑo�d����O6'��#��c}D�4�㰌�Vb�vG5#�O狮��]��ߘ���o�j��T���2�4������`ӡ��4�N��\��uu0Z �g�wy�#WEG�Z�#ؚg����}�
{�f�P�m���^ K���)V]F{�@$K;���>*�_hʊ�"�����,jW;��-�I�T��D�l�����ɗ�^�?Կ���&�V%���j!�X �eb���s[T�	��ZhJQ����l�"د��D�\JJ��ؘRo��Ƿ�+8*��X� ~=V{� �
�Y�dI��)�FдK�i��0ŽH����.��C����̓S�����:������;�Ί�c��K�K���(�*q���B�yuhn�Ϥ�5�`'I�0�M�>8Rr�?_ɀ��
�OMZ�����$���УQ��@�npB�4����l#����{�5<U��@��{o��]�������0��ӯ@�tHM(u''C�϶
Y�ߧ�~ǲ���,��"ۋ�z���������_�\k��/ɫ_�S��U�h,�����n'Hgw=�Z����������B�I�ZY��[|�lm�03X��GEH���K�Kp��Nl�-����,Bv0���ZNKS��M'cLٔ������|��e�b�7
�V��ܛ�,��8�yH�7��7w���%�ʒ�PsƓ\���R�t�'�Yp�&u�B�Xg����B`T���hM��)nC]�rm�W��y�~��$],
nJ��q�6�D�W/N�t�!��bl�u��1���c+��L���:,T�/�@�����ϱ�B`uS���%�4�k���iH��^�nIߏҲЀF��sf:Ɨ	W����>�֭�Bl8�m�6'�Y7�(�Fv�.��X)�]<�3q/���E�/�h0�ֹ��]�g��E���{j���O�h���"��Spz�w$�j�ab�jPE�k^��'R�p~��K=�߬3�J+��l�i�0W��TK�g��&=�7 C=:4��VJZ�M�@BLwFKo����@� �Y�W�cQ�*xE��0�^�ƴk��!H�?v _���ED��P/��E�����~�NI�'��\��r�s>�N�sȟ[�U��6�����h԰����f� ��'�T���*�C��e����"���̊�Q�A�!����*�bG�2��>�[P,��M�m(	�o�^S� uY��L���d������m�>�����`N�mlґni|&Rݝ�lT�`�k��	�2�S�<��L���'q�#D���I�գ@+�a�n�����pI��W��H*^�+�x�3	Rnǉ�%�1�xѴOjMȀ)ɢu��ɮ�OF�/_`������Cz&�A�n^��5{�R.t����FR��[�|GC��o����h��2�M�Ad$)�X�T���Q�M�#����Xr}� !���TYP�ޥ�Z4��/pk��pwb/hz�����R�U��	6���f')VJ�p�!i��2X4o��F�w,���z�nk��Ǿv�� �M/hW�Hk; QelՐת������um�|����8C�l�m�3��,�k��K;�����]�خ�GUFX�8�4&�ݎ����'���8����Qx��B�*p5SX�X�L�Tb����Hp�y��(�<u7q��������
��M���R6jY�"�ޭ���f�7�n���)�k�B1���:4���n�J.�G��Am��gW4g/�_�6�W��~��L�N�=�Y��iN�u�㊉gZ���� c�����ei�F/\�<����.���Qg'�>A�]6M�Xr�0%�8hb7���2�+p�ڮߥ�'z�!�>Y7��d�����$�:�΂�6d��|1@yRR��?i
 �M�K�B@ U(,V<6�k�ST �*�y�{y�(�5�<P���Y^�!�)J�"��v���h�	�-�	ȅZ�J���XvoK9����OBt�MO,@K�<����Ҋ/���߳s�"�+��&�dk�>�#�v�Dk����t�e�,��iqb��%(�ڷ�1[���=���:[�u5o�{��cd��?�Thwe�`�o,D�^.%�3�d=b|fo���g>��-_���mdKhh����{�.����w�.�=)����t,��fϡ|���@W
I��{�h��X����$<w����x~�gLtrYg7�0��D�2�t��y��R�u�!=;�
�Aui�-0����8�r���2���S������M<�+KN� /w�'�kF�Ahƛ�&�Vm�[<�۷-8C�n8�7�?=5��S*���|g��?����0lb�z���9�1��#���nr�㥏t
�!�W��W.��A@J��l�ɺݺ�����[��``���3�/?|��^s��<�hT���s>�� �����i�؛)r� sbW�p�N�W�6Zel	/0�O�4t�a_����ZC�~��!���X=g�/FC�+�g���x!�@<����1>��n�N��b"�bm�t���sB{L�'�[3��"�-��O�8���z���.ɭ�ㅭ����-(������/�؈#>����{��yK�����,�D+т�_m�C�ՑT���ᩤ�B1�V}b�S�HgL!ETt�P]�3���|�	�T�M�L;(aiY�zG�<�׀ۋm�;!ԨE5�(04 �B�TEB�;�� 2P,���1>���,<�-��F0+�]���:�w�8����p��xUg߬��1A���A24�r�H@\�����)��z�δ Q�rbe�4���3]�=z�n��Z�-�NH����!F�5��pv!��Fx�7�{��j@��V��y�<kL�0���e�q$:-Rfh�w·�l���A���C���@��s��C�i���G��&�b\��]��a�#����M,�_"@��!x���1�L,�Heי�^"Ŵos�����A��b�N'��vO����	;��M��D9z���9��������jF�q󻖔TG��(�㈆��a.�1��Ut3�T�n�m��G�L����|�A[�8gk�o�ۡG�5�*�"�:wF=���d��}|x4, e%�yo#�p�zPR���B#BMw�!��I�p��rC��`l{�����Z/���m��}Q��dNH�(��[��1��s�,	ֺ1Zu���ި�st縉��|z��4�����ʭ�A�[��ܭ*v���`��$=���*�!��wf�>��q�~7H9�1]0����n�}�W�ߚ��ֵz�R�rx�=�9K�(���
�/#NU�#�.��mF�A��Ąȗ�Bp��\d��$��55R�3��/��>(vʲ��_KK�2���5��cw�����+���R��͋�C��?J�u����#xU@���E�Z��Tԓ�y������� 8��	Z� ���~�s,�b|�ǩ ��Ssqn�O+|�������.�9?�Q?�L�Zl��؜�Y�j�:�ūƷg�sT؉*�5 �6*ͷ7�h�qL�|r����9��  0��j/�����&-��/�Ҧ���,v�\+}2�/�[������ѻH�ɷ�u����)N��v���tY�Ժ�cW��&`�A7��U��g��8���G�hǭ���2+*�$�[�f���H�%Z��U ��v�� E�A��)<�3~PKvw�orRi<�(���U���	�r$��5{�^}�9��>����.����a�	��T2ݯ��ć��햿������i���NL;�6�#1�W�ٰ��Gs�L$%Ї)�������i��NC%����,���&����x��	/��G��>�<g���Za��� v�5�hAe=?(���K�31({ B�Sˇ����<�F�z�7
4�]�q5�au����R�TZ
���+�FB��c�,�\�RT�i��?��jϼ1Q���L�Dыc�m��p������oSFa��|�>փ2�2�ǅ�_"��c�K����jR��ķM�*,v�|:7(P��t��Lk4'��H��m�'��&]]��ڲ?amm���NM��b�5�v7\�!��n�cX�e�Q���y)���Ӧn����'7��#G��W��/'�d�V9��+�m�7>-�d�V����X�T-2�n��P̅!Ӝ`:��>��e!�_퀎�GY�E�i���	�g�#������<�rM�|�e�ܽ�ѭ� �,��-
܇JVH��њ!}p������S��}d��{��:�����Z�5-�
��/j�V�w_E������tC1�ybW{1&&��K07����5�� �~H�����t�9B�� ���!���J��fdD��ʭ����)w��v��Jfr�����(Hc���ٺ��z�;q�yF�1&��$�bn?E�W�e+ȓu���>�s���Y�EeV��d����b|Ӕ�"��$t���@�1��TF4�B1s�/�SE�W��������k�bv��32�{z*���q���t:�n��+ഉf$��Qa�?C}�%>8�����M3��EP���9ʊ�Q����D��lV#��~3�W��vя$�O\��n2���,z�)�L��v	]Q�J5❗�f]O�XfN�i؅1��9���/^���s�I��l�a!�
gt�Ǖ��<(�d�����yX�Ū���b��I�� ��9�v���
mbP�t(]7�$��糐#%��������#6�뢀7E�E�g���[��ў���]�u<�F���E��=�5�a%��w���b6g�I�T���4�ʄ��~�
&^���Z�և�M�T*vި##��3ef���냼���洅�7I���ut�l��W=��0Z]iŀ`�}����x��j�u<�������_p)�� [5�dP/*����s�!�-{����.�SoD��Q2��7�F���\�}���gXX��}���e�40$�^��U��}Ca�ﺣ�-m���P�0��#�/r�L
����&;���`l�b�2S�Qv�AuWZ�28��_*���+�w��a�:�]v�A�̨�"�=ضR�G�>��e�?��'�`�A&���{��(m ����İb���;T����t�jeܐ�U���גeʧ�9��]!�dHka�UI1��(���+Y�T�X/Z��x��|�x�+��3l��7:s.5�1��
���t��>�}8[�|X��5[�qY,E�h�Qm�X��Nܰ҅���qi���(k[�ڇ��n��VK�����Z��>)rg}p`_R0p�Kb�Oɱè~��v����H������z�W_u����0���]C���	���c!����i�جq�_{��έd�H����`�8{v�6��K^+͂|
Ͻd ^AR�ƒ��e� xk�sw�F��Rf���I�?j��L<�s0F�x�Tu�U���h~2�yS�)H)@b��sO {�1����=�{j�>a���"���CG��3�/�{����c\�	z�-�0puh�0���o	�%�v ?�) ya�k��S�ݻ�(�K��LP0}���Гw�a��12O��p&H81E[��/�9rr!��(��&-h�����o�vI��>.�������@�Vn�F0i��-�܋����K�<m��&!n�ḋ1լ8��_ZbS��v[�Lr\<�(�"���I-T�H&�� �I(*-��#w�2����k��(;,���*��%���TVK�o�لC��J����\��h�&��h������4��u:@b}R\�����/�L���Q:�4�A-+Lq���Ed�X���l�{D�������,��+�ۥy��\���F�l�e�o)Yb���*�5!�$�nP�5�_R�ACۡv�m�S	F� ̨V�&z�5�Z�@M�䟄T�]�V�v�Ce��0�p�o�E�X��\�*a�T@�����/�QZ��]e�\�1��)u��ﮙ�)C���&FO�:)����,�ZX�ժ=r�����[�ݥ��6��tI�~4Q�9Y��I�ŞUe��P��1l&DQc��;�&I5��\X	�
���	��b&�ed7M5�S���4]nM�E��b\Ԓ�Ǧ� .���5���vFD;�����҂U�Flx�N�Hj��A�����z��syODPo���1a����k�C;��ٝ"$�c	�W�U�O7���F���}6~���XK�1��í ��`/��2cAqsD_ R�;;���6��\p_U|��9�5^%��c1���j:��3�X�t�޶�D��L�_�T/�B�,Oyq�u�w���4:�r�&1ץ�!	�����z���Ō�3.Q�I>,�r�Uݎ�C~)���5�L�Ī����d=����mn�1B�] �4��ĳ� ��DErk[0���I�C����%s��Xޒ�,{��
ʞl���9(�����m��(�: 5Z����A��}$u~PG8�1� ҟ�(����&{Բ{�2��"�'�p�ց��:k��nMy5$�� 7U�>�FNf��0d�'�a:����>���c#ȶi�(�E�?\�.xIo���&��� I\4~�f��������t���\zy��j�^zf�^����#)eW�0�j ���[�.\�6G�I!,���(*�5���o��	���*0��_B�,�^%��b��DI�	��� c8dH�`U`kos��[�"~i�WZȽ��I<j3ۓ�N�.�j�<�p��+��&�}o����������у��)��@�$�C=�.(�[��=�x{m�;����?������N�TϑpW��(��lܯ�=?]z�.ƚm(����ǒp7��˩"Z��ksN�6ۖ�'��K�]�ؼa��g�Q�w�����i��xK����F�c1.�Ob�@��87�J��O�*���G.�U��oC�����ԟ�d&�O��:Ow��ߑ7�Hd���_	�_$n�P��p��*\B�dڹ�?�wbzŴ����g���9�ϑ�O��J�mc�N���C�d;���?���|�O�� �Z���jw2�k��@�hm��"�.N�V��<r��xۤ+@���)c�찁��/-9n���!�� Z;7Bx.��O�Lr?�v���@��x��=����i^5�/l�G���7K�,X�O,w��zg�� O�$��hDgNM��	�9���_�cz͟��ӁH�{bu|�=�I��!�FS8F��98�Oq�;�=TP�[:FX�_��ŏv��Ɵ���w���B2��!����OeX���m!v��<�A`��Z�8«]���.�x���ɈX#m�6m�����v����t�8'���r�rU���n[�v�ӆ�gh���G�dx�"��c�,B
p�c�bN�K�l>�?����5�R�k�N����W���h�'\����F��J�݋:E&Z��Щ����|t܅�S����^nZ»�}���4,cnݑ4�G=d� ���!�1"́ܥF���U�Ȗ%���ц-b�\q��w�Tnbǎ}/o��D[�D
�fT�r�BJ�����n��g'��f����W��Ti���U��3?��b� s�7.������p��W�������,%8��CfZ4�@��w)8�=Tr��9�����{��I�_�K)|�������Z��N�`�m�3R���D_/���(����u��R���?s7�E��*s�-��:�� ɗ�z95	��Jvw"�\��/�B�è�����:*�Y�8|��?������x#��ӳ�ZmW�|k0��dc�@����Z5�x��аZ�*��� VU���g�z���$�:+"��au�\V�����-[��U�J� ����o��pٔp�l��+�M��qH�\������5�f��Z�U�Q�v�ƨ@�xQ�T/qS@֧]�5��v��$����=�H��D���9"	a5O��c��Q>�~լ��J����M����(��>?�ٕ��P�h���7���[6�S�z%�42�2�Qi�m�]�߀D����J'�ˎG�ѧ@��r�5I�Y��E<�s��u��N6S�� q g�N?BS�v}vYl�Ũ�&C>�,�Z�{W�,���In����C�P|`$ҙ\���!j���*54=e9�#�d��w�ש�	��Q�k�>��������+x����C� a�Ql��h�_H|ֺsQɸ�d�J�"��HƘ/%!o� b,�_#��`�w�����\�j:�t�j)��j�ql���U[k�� [����#q�'��b��WݲX3wY��c�l�C*��P>$�;Z�4���d�� S$
�]�Wqr9s�ս�$������7��@��;,/hR;����0��t�"�gM�ı��d����1*U��bf��)������vU���.8Dx�N��B�D?�����V��C{���~j�L���2@�|{SP��#��Kڰ���ȏ9L���b�����Ɇ�"��[�Wa�
F�]/9�p/�!�Ϸ���H�zx$��!�LF[�y�+�儫[�����ǜ�f�?���������]���T�e-�
q:!1#;$�ؙ|����Z-�n틅���S�˳]��B9�����
���%���=,!���X�~��ĦLӊY;�#��0�(o� �D��2Ԓ�M'#�
Q���>�3�6��=�� n�7L�W�.uv!���M&7��,	�'����ܥ��y����֭(��o��V%J�፯�ɶ[��؇��臊��JE�w�SR���-�!t��i]7
aM���]Q#¦��~�(�~㶔=HH�N8)�2n��2ؽ�4����i��U����@���;���Q�$�� qx�a	ه�3k��N��=3N��O}N��%Q�tJ�s��Z�YlN�Q��5����fa�|����r�␰��xc�h+��%b�hb�=60�T*~woބ�4�.��ofrD��u�����sz3w�F��=eӑ�|ኩ�������4}���M.iv���6�_�P��bb]����G���F�����Wgs�Q>4?��U�t�����T��h�L�����ك~.	4��R�È��=H�A�ԅau;���������<�Y��ӅE,p�SU-�X4 8 L��y���l�w�7ګ�!	~�*�&,9���U�;��!�_txإn�L"]�`��<����	Ƶ"f��+��K8#g&�Ĉ��:�mB������:I<ך
JË�j �d5v�F��]� W`�v�:s�b����X��}T���z�����<-WA��N�-�Qᗨ~+=���g\��o����Z�#M�௳Z��&����N� x�Gd���й��{N7�ueY~���7՜4�ZN� z�A������.X��A���j\Uh&AuX�8D��}Q~i5%�^C�Kx�c`&��N�	}w���,Dw��R^�Ne�x��n���|�Bt������eV�iF�D�Ҙ_Cm�Nc!b���h�g�)�����#BAUy�D?P?�xƸY�F�^�9Ho��\p� �L��$��"6<���"uِ^Аgy:z��8�g�<�^��lLP#�Y�
⢑R�fP�JC6�$��qІx&��.�t܍������c��Y"S�� zS�Zl�(Z���0�~�SE����­ #&���࢛��ezj�yY��4�0c��i��������D���(��j�8Ș� �qtD��%-��W9����N����*��ax9�f�$U��	��/+2�Da��$3?�O�ƫ�-��>K<��M�^��N|�Y}�TK�U���~�Ag�a�A�炪t8���G�t�T���.���}��\�(7�١��J����8rQՋA]�/��
�E�.B��X�Զ�2Wg��-ć�~� �:�範v"a�	ϤvC�CIl���T���Y+��/�]�㈷��=�����2��+_t)F]�f��f��7K
�d��o�v���lh;ۚ�f,c%�qiy�=���{�5)G*�M��/�VHa�nƬI>�
%uTٗ~�>���`�+�`G�_3v���Yzz'��UĊ�v�9[���
`Γ^��H�q�<��̓b�|Q����i�o�w �6ӵ��Ld�� �#ʌ���eY��U'�|�h�^�8����׶O��F��Ԁ>���U����`���Փ0ܒ�{BCR�/.�6��C{���\,W3��)����Z�|��b�֩r��V|ir�l	P���Ӆ��|�Ck�����J����m�"�j���8���@� y��B����Y�R���e/B�*vMg��ƐH� {Tg��;��˨��5I�\M��h^KW�ƃ��`�Z�%5ћV��ha5�,ԏ��ک�����ʢ���1��v:!�	�Z �?q��=0����j��4_!�+o���q?�'%Zg]�JBJ��L�¥����P����z�/a{{�K�M�D���V
$�Tj��w��\����kv���,{Ŧ��la�G�I_M+F|���V� �b1XR��9�0�P�/��0aRʳ��K���a��&.\l��}��>��,�F]Y�gT3'��+P߮�a^��*8G#��s�/��@���L-b�X�{]?�ȕ���[?�P�42|��y<�(Yg�7ǀ���m�\���r����[�lK8�6�Hxr��0l�_co��ȇ!.�{��՟٦2饿�mT6|H�6b�
$ӾӋ����,ёZ���B�`��℆�#�7�]B5�4�